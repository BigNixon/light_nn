package my_package;

    integer connection [985:0];

    localparam integer network_structure [3:0] = '{10, 64, 128, 784};  //     10,64,128,28x28  
    localparam integer connectionRange [4:0] = '{986,976,912,784,0};   //    ans+10 , ans+64, ans+128, 28x28=784, 0
    localparam integer weigths [109385:0] = '{-53, -114, 105, 172, -122, -190, -238, -76, 123, 128, 174, -250, 101, 76, -28, 186, 93, -151, 84, 136, 122, 150, -222, -11, 137, -13, -137, -155, 229, -138, 43, 153, 85, 130, -30, -176, -10, 56, 94, 64, 119, -102, -134, -203, 141, 17, -177, 4, 4, -195, -49, -192, 35, 0, -26, 92, -139, -182, -83, -171, 122, -144, -164, -60, -34, -259, -195, -56, -184, 87, 35, 123, -35, 22, 67, -216, 119, -177, -125, -157, -89, -66, -182, 37, 61, 102, 43, -163, 203, -62, 39, 47, -21, 168, 147, 63, 124, 115, -31, -70, -48, 67, 21, 147, -200, 117, -194, -33, 136, -4, -262, 48, 65, -118, 73, 151, -51, -116, -171, -33, -207, 146, -123, -127, 51, 101, -204, 117, 95, -221, 241, 169, 46, -218, -238, 8, 117, 126, 19, 126, -89, -86, 133, 115, 188, 64, 123, -56, -189, 27, 134, -89, 122, -212, -35, 113, -58, -121, -197, 168, 28, -289, -30, 106, 170, -71, 101, 35, 32, 138, -233, -54, -129, -92, -207, 7, -190, 129, -151, 17, -219, -128, 54, -112, 169, -48, -211, 188, -86, -116, -93, 46, -99, -271, 149, -656, -166, -30, 145, 22, -108, -216, -112, 63, -104, -267, 62, -134, -260, -181, 101, 69, 105, 120, -319, -248, 103, 37, 136, 30, -179, 45, -157, -34, -122, -181, -124, 46, -287, -206, -190, -30, -102, -172, 38, -157, -188, 160, -62, -141, 92, 78, -231, 193, 52, 124, 188, 147, -105, 133, 93, 165, 63, 49, 168, 140, 52, 114, 21, 13, 23, 139, -136, -32, 56, -169, -86, 180, 23, -132, -113, 49, 144, -150, 33, 75, -196, 192, 38, -66, -213, 101, 93, -197, 148, 130, 50, -168, -13, 96, -277, 75, -248, -23, -144, 144, 133, -152, 11, -142, 53, 33, 26, 33, 84, 63, 83, -227, -207, -1, 125, -225, 66, -150, 11, 160, 26, -174, 125, -219, 49, 43, 108, 92, -79, -10, -141, -282, 118, -154, 188, -80, -165, -174, -170, 183, 58, -167, 90, -40, -206, 153, 140, 107, -34, 51, -25, 98, -118, 117, 95, 156, -37, -212, 10, 34, -69, 106, 63, -15, -175, 18, -48, 64, 46, -92, -49, -72, -241, 122, 154, 50, 84, -99, -243, 20, 144, 11, 198, -76, -79, -154, -88, 37, 140, 25, -211, 29, -232, -17, 188, -166, 120, -148, 43, 163, 102, 163, 50, -47, -136, -121, 117, 158, 27, -99, -141, -18, -255, 94, -48, -113, 173, -35, -197, 102, -206, 15, -109, -62, 111, 173, 55, 92, -138, 38, 133, 125, -181, -147, 10, 49, -140, -52, 154, 108, 57, -159, -141, 175, -202, -144, 99, -169, -87, -142, 144, -7, -111, -39, -209, 92, -150, 80, -85, -14, -46, 43, -26, -75, 30, 138, -179, -144, 5, -4, 106, 88, 120, -176, -47, -53, -109, -160, 52, 39, -150, 112, 145, -227, -131, 73, 141, -45, 27, -85, -108, 84, -189, 185, 180, -190, 114, -79, 4, -75, 185, 188, -105, -215, -32, 2, 27, 197, 116, -18, 78, -268, 39, 1, 71, -199, 144, -121, 80, -163, -91, -172, 132, 189, 1183, -16, 98, 72, 165, 58, 139, -189, 108, -151, -47, -157, 144, -164, 168, -82, -189, -55, -196, -238, -147, -211, -77, 17, -149, 103, 63, 142, -35, -124, 150, -184, 145, -171, -125, 17, 20, 97, -103, 125, 96, -57, 94, 124, 39, -176, 91, 88, -48, -162, 42, -187, -119, 120, 184, 146, -112, 143, 174, -118, 55, -132, -170, -175, -122, -869, 156, 43, -173, 30, -103, -39, 77, -8, 134, 66, 96, -202, 92, 68, 104, 9, 101, 154, 13, -105, 14, -54, 39, 110, -263, -152, 78, 129, -216, -135, 96, -131, -185, 156, -114, -245, -225, 35, -56, 57, 58, -137, 111, -266, -84, -251, -186, 173, -139, -192, 157, 90, 129, -34, 71, 42, 105, 6, 97, -218, 59, 15, 46, -154, -48, -23, -37, 8, 143, 18, -66, -10, 12, -15, -69, 26, -70, 66, -23, 59, -24, 118, 76, 31, 1, -30, -134, 108, 85, -49, 79, 256, 4, -108, 8, -35, -23, -5, 29, -133, 8, 5, 54, 29, -11, -24, 10, 164, -33, 20, 84, 54, 65, 63, -82, 45, 104, -31, 42, 94, -32, 5, 108, 40, 6, 11, -55, 95, 36, 67, -53, 98, -4, 10, -12, 151, -135, -154, 145, -63, 85, 35, 93, 12, 25, 105, 49, 149, -56, -26, 86, -12, 71, -38, -32, 45, 32, -77, 45, -45, -18, -46, -40, 82, 105, 46, 6, 31, -71, 66, 45, 11, -14, -7, 32, -32, 48, -80, -15, -69, -131, 41, -86, 13, 58, -136, 50, -128, -52, -90, -97, -52, -112, 202, -44, 28, 87, -8, -124, 23, -86, -83, -58, -2, 66, 47, 65, -19, 14, 84, 51, -95, -39, -122, -32, 80, 22, -43, -10, -76, 110, 58, 107, -15, 7, 22, 54, -10, 17, 84, 136, 85, 77, -91, 13, 5, -111, 24, -90, -101, 60, -107, 52, -32, -27, 90, 53, 42, 114, -23, -69, -3, 50, 136, -96, -52, -116, 44, -87, 43, -19, 29, -12, -106, -23, -24, 79, -22, 69, 78, 28, 10, 113, 40, 65, -73, -132, 70, -76, -42, 60, -74, -65, 168, 122, 142, -11, 111, 4, -44, -17, -38, -4, -158, 49, -8, -86, -10, -58, 122, 177, 82, 40, -144, -58, 67, 12, 31, -120, -24, -59, 4, 60, -70, -13, -51, 107, 60, 62, 25, 35, 14, 127, 46, -63, 32, -19, -144, -87, 37, 33, -81, -95, -146, 1, -105, 107, 0, 127, -94, 43, -91, 67, -12, -2, -28, -82, -39, 6, -255, -1, -30, 24, 45, -33, 109, 19, 76, -29, 58, -100, -40, -3, 54, 128, 24, 21, 44, 104, -162, 97, 2, -36, -100, -108, 160, -31, -176, 39, 48, 37, -47, 13, 18, 66, 99, -1, 125, -8, 51, -101, -37, 115, -121, 41, -59, 183, -96, -56, 154, 250, -88, 114, 32, 38, -12, -78, 58, 2, 20, -21, 16, -47, -126, -2, 76, -25, 101, -67, 13, 3, -129, 28, -130, -56, 35, 92, -23, -21, 19, -50, 12, -17, -52, 94, -12, 60, 11, 12, -103, 57, -54, -129, 94, 4, 20, 113, 60, -94, 166, 158, 260, 75, -29, -92, 118, 60, 4, -18, 92, 103, 62, -38, -65, 18, 15, -136, -39, 59, 98, 12, -82, -30, 19, 82, 116, -83, 17, -86, 63, -12, 46, 73, 103, -97, -28, 28, 11, 35, 73, -6, -32, 59, -88, -89, 35, 14, 97, 8, -118, 11, -50, 118, -53, -16, -70, -36, -109, 18, -14, 56, 57, -59, -5, 55, 13, 48, -35, -138, 48, -27, -61, 81, 55, 14, 138, 95, 32, -97, 96, 73, -59, -23, 48, -122, -50, 140, -120, -55, 90, -92, -30, 12, -67, -119, -4, -71, 106, -49, 71, 39, 0, 52, 56, -15, -6, 55, -101, -12, 20, -76, 1, 90, -17, 2, -109, -14, -39, 63, 10, -57, 65, -36, -8, -11, 3, -47, 37, -33, -11, -188, 43, -10, -33, -24, 176, 43, 31, 1, 172, 85, 149, 61, -115, -53, -23, -79, 27, 0, -30, -33, 39, 229, -138, 18, -3, -31, -5, -80, 106, -34, 21, -9, 3, 31, -9, 28, -76, -34, -19, 218, 40, -9, -84, 15, 13, -115, -28, 78, -45, 58, 36, 16, 13, -2, 66, 65, 93, -18, -86, -47, 28, -16, -174, 37, -153, 16, 77, 49, -36, 126, 9, 29, 180, -93, -29, -259, -82, 54, 5, 20, -166, -10, 76, 84, 18, 3, -84, -111, 116, -24, 44, -21, 3, -149, -51, 30, -33, -87, 19, -93, 5, -140, 28, -7, 56, -114, -25, -83, 31, 22, -9, 11, 27, -58, 65, 79, 8, -8, -70, 18, 39, -42, -25, 59, -92, -2, -63, 23, -300, -50, 31, -20, -94, 247, 138, -29, 37, 74, 92, 247, 18, 13, -56, -67, 36, -1, -13, 81, -12, 110, 159, -49, 104, 110, -56, 154, -27, 68, 7, -5, 41, -86, -108, -15, 40, 38, -61, 7, 139, -98, -57, -76, 9, -93, -87, 67, -176, -103, 31, -48, 145, -78, 54, 183, -32, -46, -1, -66, 21, -4, -125, -178, 114, -199, -53, 29, 41, 26, -6, 41, -72, 146, 11, 23, 1, -160, 3, 81, -136, 13, -75, -65, 86, -106, 6, -52, -30, 27, 33, 185, 67, -34, -4, 84, 24, 23, 52, 0, -59, 89, -72, 47, -23, 37, -51, 68, 17, 3, -7, -8, -67, 6, -94, -54, 9, -27, 17, 6, 76, -57, -28, 56, -37, -1, 46, -34, -67, -142, 55, 27, -52, 196, -160, 79, 34, -99, -15, -44, 38, 14, 12, -143, 94, -166, 109, 3, 102, -57, 0, -15, 115, 76, -56, -6, 203, -54, -49, 46, 17, 33, 84, 108, -130, 60, -63, 26, 6, -39, -65, 25, 103, -29, 37, -62, 111, 73, 45, 70, 2, 19, -114, -33, -30, -128, -10, -43, 78, 123, 67, -10, 86, -58, 45, 72, -19, 67, -16, -69, 129, 8, 5, 5, 83, 135, -95, -85, 39, -30, -28, 61, 28, -43, 81, -4, -56, -66, -114, 39, 142, -35, -121, -19, -116, 49, -46, -37, 96, -65, 77, 15, -11, -24, 97, 0, -43, 65, -87, -50, 29, -71, -75, -101, 4, -125, 43, -40, -40, 33, -26, 12, -73, -10, -121, 5, -232, -39, -42, 4, 12, 23, 100, -140, 17, -26, -15, -73, 11, -70, -20, -72, 22, -45, 8, -42, -16, 42, -87, -15, -33, 231, -8, -53, -46, -49, 10, -28, 90, 71, -6, 7, 114, 46, 57, 46, 57, 112, -108, -41, -1, -18, 62, -43, 126, -56, -18, 61, 18, 16, -105, 109, -19, -83, -29, -84, 29, 68, 140, -26, -19, 207, -72, 167, 108, -74, -34, -46, -115, 7, 40, -56, 205, 22, 154, 105, 148, -52, 38, -62, -4, -113, -47, 75, -38, 69, 40, -118, 106, 18, -27, -66, 104, -13, 39, -71, 36, 11, -20, -33, 64, -67, 5, -53, 63, 48, 56, -54, -106, -9, 12, -45, -61, -55, -21, -4, 12, -19, -30, 41, 23, 53, 17, -10, -14, 17, 48, 121, -117, -79, 70, -97, -17, -28, -119, -155, -86, 10, -75, 25, 78, -15, 47, -95, -25, -111, 1, 31, 6, -66, -35, 59, 32, 25, 198, 58, 27, 1, -194, 33, 4, -5, 1, 49, 72, 2, 55, -226, -78, 19, -69, 45, -83, -72, -15, -102, -45, 43, -29, 15, -1, 40, -88, 34, -170, -35, 37, 37, -24, -61, -87, -117, -57, -10, -39, -43, 81, -208, -31, -10, -11, -194, 1, 133, 45, -117, 97, -40, 107, -18, -95, 61, -19, -10, 46, 44, -117, 11, -80, 63, -44, 30, -141, 31, -19, -4, 71, -50, 66, 37, -114, 36, -8, 139, 114, 65, 22, -92, 2, 61, 62, 21, -79, -8, -107, 41, 154, 74, 2, 15, 65, -28, -12, 75, -14, -98, 50, -104, -133, 10, -31, -192, -158, 54, -64, -127, -89, -103, 26, -29, 19, 90, -29, -31, 59, -89, -8, 29, -1, -161, -95, 21, 61, -174, 16, 3, -49, 100, -24, 68, 23, -30, -21, 9, -6, 38, 38, 42, 72, -4, 59, 24, 74, -122, 174, 72, -20, -18, -218, 129, -34, -200, 110, 72, -80, 50, -79, -12, 74, -178, -86, -99, 4, 91, -13, 3, 93, -61, 1, -74, 47, -48, 8, 210, 58, 31, 70, 27, -15, 54, 53, 37, 87, 68, -94, 27, -222, -125, -96, 39, -185, 6, -79, 21, -82, -24, 17, -9, -95, -35, 29, -22, -82, -21, -21, 64, 54, -104, 132, -33, 68, -27, 74, -66, 31, -23, -2, 5, -19, -27, 108, -65, -103, 188, 51, 297, 73, 53, -14, -95, 168, 63, 77, -91, 70, -3, -25, 48, 53, 34, -65, 54, -83, -133, -14, 10, -7, -95, -93, 24, 82, 4, 122, 27, -112, -58, -148, -42, -144, -80, 13, -78, -49, 21, -88, -34, 141, -112, 60, -90, 104, -1, 31, -62, -173, -31, 88, 27, -133, 57, -46, -19, 78, -68, -8, -160, 55, -1, -76, -34, -37, -142, -19, -13, 10, 97, 59, 42, -38, -179, 26, 7, -164, -154, 98, -43, 19, 92, 79, -92, 13, -15, -32, 128, 62, 1, -93, -41, -56, -1, 5, 8, 48, 37, 19, 76, 70, 97, 127, 137, 2, -58, -123, -60, -49, 103, -12, 3, 97, 19, 106, 17, 176, -59, -36, 80, -27, -36, -32, -58, 11, 69, -100, -43, -157, -39, 84, 44, 193, -60, 42, -3, 61, 4, -16, 128, -23, 2, -49, 137, 99, 181, 187, 27, 19, 75, -8, 198, 43, -34, -57, -63, -16, 17, 13, 225, 33, 132, 87, -56, 50, 64, 19, 67, -30, -152, 34, -17, -16, -40, -39, 150, 38, 204, -16, -8, 122, -20, 19, 198, -21, -114, 32, -13, 102, -17, -94, 90, 204, 56, 23, 8, 36, -43, -13, 44, -20, 34, 157, -12, 119, 57, 59, -123, 20, -11, 66, 66, 20, -39, 76, -51, -166, 38, 100, 175, 150, 36, -13, 76, -10, -100, -16, -36, -54, -50, -11, -46, -114, -46, 35, 120, 87, 51, -89, -37, 17, -87, 48, -86, -25, -56, -62, -24, 56, -85, -5, -23, -83, 91, -65, 7, 44, -8, -77, -16, 92, -1, -95, -23, -7, -134, -55, 10, 179, 75, 17, -25, 152, -62, 42, -47, -65, -65, 2, 95, -148, 7, -14, -51, 26, 30, 156, -29, 42, -31, 129, -4, -73, 8, 86, 2, 23, 100, -24, 49, -21, 12, -61, -190, 30, 60, 18, 57, -10, 85, -57, 12, 18, 128, 54, -80, 37, -30, 57, 23, -233, 32, -178, 79, 147, 19, 52, 38, -36, -59, 102, -211, -34, -36, 70, -198, 74, 71, 80, -60, 155, 161, -42, 126, 26, -134, 47, -79, 13, 72, 96, -152, -55, -23, 49, -61, 76, -136, 10, -109, 16, 15, 29, 71, 72, 22, 80, -49, -19, 70, -13, 111, -49, 14, -34, -64, 86, 35, -98, -85, 4, 17, -24, 35, 30, -33, -134, 34, 44, 26, 62, -28, -4, -53, 73, 38, 0, 85, -55, 6, -41, 107, -135, 183, 64, 56, -96, 28, 65, 78, 98, -28, -1, 236, -66, 53, 4, 99, 26, 104, 81, -103, 55, -26, 139, 91, 36, -7, 94, 181, 12, -27, 59, 100, 153, 162, 13, 8, -26, 121, -1, -17, 61, -34, 67, -26, 124, -6, -90, 64, 49, -21, 1, 97, 95, 5, 36, 114, -80, -63, 219, -51, 43, 88, 154, 52, 91, 34, -53, -3, 66, 5, 30, -21, 8, -51, 85, 67, -33, -55, 65, -27, 6, -92, -111, 62, -46, -24, -101, -66, -86, 53, 25, -45, 36, -39, 46, 16, 44, -120, -80, 3, -108, 22, -55, -3, 46, -55, -35, -17, -3, -56, -78, 18, -71, 117, -65, -8, 87, 85, -208, -110, -63, -53, -174, -90, -149, 6, 88, 36, -16, 74, 61, -14, 33, 40, -15, -162, 131, -65, -83, 20, 78, 53, -69, -41, -27, -36, 40, 21, -2, 43, 100, 37, 86, -216, 10, 35, 105, 37, -24, 18, 38, 7, 85, -4, -59, 45, 26, 11, -49, 10, -73, 56, 49, 49, -28, 8, 186, -95, 150, -7, 2, -13, 20, -144, 5, 4, -225, -100, 15, 234, 132, -106, -63, 30, 126, 56, -93, -95, 9, -33, 100, 82, -126, 90, -59, 19, 22, 110, -6, -48, 2, 29, 21, 58, 22, 93, 6, -37, -29, 159, 91, 39, 16, -119, -33, 12, 4, 16, -76, -15, -78, -44, 59, 12, -27, 3, 8, 25, 6, 4, -12, -48, -45, -20, -49, 101, -203, -3, -98, 33, -28, -93, -45, -56, 71, 33, -45, 93, -33, -90, -136, -25, 48, -37, 28, -93, -89, 38, 13, 151, 23, 38, -40, -94, -106, 90, 39, 43, -54, -21, -1, 26, -11, 103, 48, 57, 50, 92, -52, -34, 100, -61, 71, -81, -15, 30, 0, -10, 152, 18, 79, -21, -74, 30, 31, 11, -120, 33, 24, 93, -43, 49, -25, -121, 19, -102, -200, -10, -135, 121, -105, -21, 121, 35, 19, 47, -10, -49, -47, 58, 52, 71, 101, -119, 8, 159, 117, 46, -75, 52, -112, -65, -4, -12, -89, 21, 66, -1, 113, -91, -59, 21, -18, -100, 2, 63, 138, 3, 45, 53, 5, -2, -94, 0, -56, -21, 36, -2, -35, 40, -17, 99, 150, 26, 51, 122, -95, -47, 80, 60, 84, -112, -129, 19, -20, 13, 66, -49, 88, 95, -62, -2, -70, -59, 37, -23, -78, 62, 81, 40, -103, -21, 67, -11, 50, 87, -56, -55, -81, 83, -76, 7, 132, 2, 182, -79, 101, 70, 95, 123, 10, -34, 57, -55, 25, -12, -43, -25, 151, 18, -20, -20, 45, 51, 172, -68, 145, -43, 51, 37, -66, 167, 140, -24, -92, 142, -21, -11, -25, 126, 11, 124, 21, 87, 166, -123, 38, 34, 34, 88, 59, -5, -77, -115, -22, 21, -1, -41, -45, 25, -2, 90, -60, -4, 120, -13, -26, -51, -174, -37, -85, 84, -14, 61, -20, -49, 105, -31, 124, -56, -89, -34, -39, -38, -110, -6, -35, -64, -60, -41, 299, -32, -63, -39, 31, -113, -108, 24, -62, -108, -33, -226, -4, -4, 102, -94, -49, -68, -48, -69, 83, -92, -137, -11, -68, -41, 94, -150, 52, -128, 18, -85, 29, -20, -4, 111, -56, -50, -47, -49, -97, 95, -33, 22, -34, 62, 77, -106, 28, 12, -32, 71, -164, 53, -100, -257, -11, 23, -41, 82, -28, 43, 109, 98, -186, 121, -45, -3, -57, 73, 4, -38, 103, -179, -22, -55, 87, 69, -58, 53, 57, 51, 72, -24, -118, 148, -17, 96, 114, -92, -81, -165, -155, -54, 31, -86, -43, 93, 69, 8, 110, -48, 36, 57, 30, 30, -6, -93, -62, -19, 75, -46, 26, 80, 49, 54, -9, 52, 123, -43, -8, 77, 7, -32, 79, -22, -93, -15, 14, 307, -164, -39, 22, 52, -113, 86, 36, -157, -128, 52, 145, 60, 6, 4, 91, -10, -72, -1, 3, 39, -6, 46, -82, -25, 25, 18, -105, 7, 85, 12, 6, 23, 65, 35, -62, 26, 3, -75, 58, -24, -19, -64, -60, 62, -100, -166, -35, -111, -19, 94, -52, 27, -36, -30, -13, -71, -22, -103, 134, -32, 23, 66, -157, -9, -99, 107, -100, -5, 71, -135, -67, 35, 111, -217, -38, 141, 44, -166, 80, -28, 100, -27, -8, 137, 16, -23, -51, -86, 18, -68, 56, 30, -6, -158, -44, 25, 59, -41, 67, -45, 117, 12, -22, 36, -48, 44, 69, 3, 62, -84, 3, 2, -15, 39, -83, 84, -75, 24, 125, 38, -39, -38, 63, -72, -62, 23, -108, -69, -5, -142, -61, 35, -174, 78, -29, -39, -77, -42, 88, 88, 102, -41, 13, 72, 24, -163, -115, -11, 106, 63, -33, -102, -15, 145, 37, 28, 36, 20, 26, -34, -12, 21, -63, 23, -21, 6, -99, 53, -5, -120, 4, -113, 96, -57, -51, -115, 10, -49, 59, -92, 76, -35, -66, 1, 94, -94, -49, -43, 29, 45, -29, -233, -4, -127, 15, 41, -15, 129, -102, -159, 7, 28, -170, -40, -6, -14, -208, -3, -44, -32, -53, 58, 110, -12, 67, 2, -97, 19, -85, -8, 59, 98, -100, -54, 8, 56, -28, 3, -25, -1, 7, -100, -24, -8, 9, 20, 50, 55, 20, -28, -21, 87, 135, -65, 105, -7, 72, 111, 8, 69, 17, 75, 16, -13, 29, -7, -18, 159, -26, 4, 2, 30, -171, -85, 73, -87, -132, -33, -219, -4, -21, 3, -32, -12, -104, -25, -2, 44, -113, -229, 45, -44, -34, 97, -158, -18, -82, 68, -2, 30, 11, 16, 34, -34, -18, -56, 44, -208, 47, 14, -8, -43, 71, 123, -63, 2, -38, -10, 50, -102, -24, -122, -114, -29, -35, -27, 72, 36, 16, 40, 175, -97, 166, -35, -101, -69, 73, -71, -18, 28, -161, -38, 38, 124, 79, -90, -84, -3, 23, 83, -54, -65, 104, -70, 78, 50, -75, -54, -58, -131, -37, 38, -62, 25, 21, 67, 4, 118, -23, 138, 8, 3, -20, 64, -41, 28, -69, -26, -26, -12, 57, -18, 38, -8, 51, 9, 75, -15, 80, 85, 6, 27, -22, -56, -28, 43, -49, 138, 89, 78, 135, 23, 98, 26, -32, 112, -13, 217, 54, -16, -28, 84, 65, 137, 40, -12, -14, -5, 41, 16, 28, 46, -56, 79, -75, -17, -51, 88, -15, 101, 1, -107, 11, -53, -65, -36, 119, -47, 11, 110, -39, 83, -99, 149, 37, 43, -44, 21, 242, -163, 120, 178, -60, 85, 57, -50, 0, -2, -45, 74, 158, -57, 19, -10, 75, -74, 159, 108, -82, 54, -146, 84, -145, -63, -88, -72, 68, -70, -30, 163, -2, -54, 47, -93, -72, 208, -1, 130, 37, 34, 0, 2, 39, 2, -19, 42, -69, -18, -29, 125, -52, 30, 22, 3, -17, 33, 19, 40, -113, -4, 53, 35, 14, 129, -124, -57, 25, -100, -104, -94, -107, -33, 35, -189, -17, 140, 21, -65, -24, -197, 147, -18, -65, -54, -10, 1, -41, 1, 15, 105, -194, 140, -92, -159, -77, -24, 16, -71, -30, -21, 13, -20, -69, 61, -36, -30, -187, 1, -185, -113, 28, -72, 21, -36, 12, -54, 19, -92, -186, -19, -74, -32, -98, -175, -169, 8, -1, -8, -25, -23, -24, 7, -9, -72, -11, -46, -46, 15, -116, -40, -65, -53, -135, -102, -12, -48, -65, 93, 78, -117, 16, 6, -119, -18, 86, -54, 59, -39, -158, 27, 23, -119, 75, 99, -49, 50, -100, 49, 16, 80, 7, 34, 72, 82, 12, 17, 72, 66, 45, 132, -91, 31, 79, -21, 45, -94, -49, 29, 87, -21, 25, 38, -29, 66, 13, 5, 7, -55, 94, 55, 80, 93, 126, 51, 168, -28, 11, 35, 43, -147, -124, 83, -29, -77, -59, -168, -62, -11, 33, 88, -46, -56, 15, -6, 29, -82, -139, 71, -19, 3, 193, 116, 7, -36, 11, -46, -9, 38, 95, -39, -5, -4, 41, 7, -75, -3, 80, 182, -63, 115, 170, -4, 121, 39, 16, 7, -141, 115, 7, -152, 41, 7, 3, 50, -38, 24, 80, 158, -108, 163, 9, 14, 9, 53, 44, 3, -6, -187, 27, -81, 70, 98, 46, -66, 60, -4, 68, 144, -85, 93, 43, 113, 70, -40, -138, -121, -129, -16, -29, -52, -75, 24, -18, -36, 116, -104, 53, -76, 31, -23, 46, -113, 22, -34, 21, -3, 97, 58, 91, 0, -103, 53, -43, 6, 16, 13, 91, -121, 32, -47, -69, -19, 24, -126, -41, -41, -88, 28, -25, 42, 43, 56, 151, 52, 18, -61, -59, -111, 104, -133, 34, 178, 121, 52, 135, 68, 98, 50, 53, 5, -26, -73, -16, 139, 138, 78, 209, 106, -46, 57, -106, -36, 11, 94, -46, 30, -3, -12, 76, 48, 66, 122, 147, 94, -55, -86, 79, -75, -48, 20, 4, 11, 17, 79, 99, -39, 82, 32, 2, -8, 22, 59, 46, -11, 4, 51, 77, 127, 39, -32, 26, 64, -150, -116, -57, 13, 117, 51, 43, 99, -115, -67, -59, -46, 139, 0, -11, -68, -93, 60, -109, -83, -10, 54, -81, -55, -98, -72, 111, -81, -106, 44, 11, 32, 61, -32, -80, 30, 79, -36, -61, -62, -76, 42, 46, 160, -50, -45, -28, -12, -146, 37, -32, 24, 87, -22, -94, 249, -15, 62, 125, 95, 30, -45, -48, 54, 24, -41, 181, -29, 115, -43, 97, 16, -59, -37, 37, 52, 45, -85, 14, -59, -24, -56, 46, -105, -108, 55, -36, -108, -83, -130, 90, 16, -23, 59, -56, 72, 112, -60, 36, -38, -41, 41, 28, 26, -63, 44, 46, 39, 58, -70, -110, 32, 40, 65, 5, 30, -146, 75, 17, -33, 149, -45, -1, -13, 92, -4, -101, -130, 132, -47, -31, 10, 36, 115, -51, -40, -1, -111, 43, 72, -83, -65, -44, 15, 62, 204, 14, 31, 18, -61, 139, -34, -14, 98, 17, 48, -99, -100, -80, -50, 140, -14, -35, 56, -23, 65, 51, 29, -39, -98, -21, 59, 55, -38, -6, 93, 5, -28, 45, -160, 11, -21, -27, 36, 118, 55, -18, 56, 85, 27, 73, -22, 48, 36, -167, 2, 54, 25, -28, -81, 42, 152, -119, -25, 33, -21, 65, 6, 115, -43, 33, -5, -126, -93, -63, 67, 28, 85, 28, 22, 37, -50, -25, 62, -122, -67, 38, -109, 61, -102, -14, 23, 35, 39, -2, -15, 7, -46, -11, -110, -28, 27, -254, 54, -137, -37, -15, 69, -107, 61, 29, 2, 160, 113, -5, -66, -80, 132, 185, -45, 44, -55, -18, 147, -20, 30, -56, 15, 12, -48, -4, 100, -7, -111, 86, 18, 62, 42, -3, -140, 101, -113, 12, 43, -52, -58, 112, 26, 64, -13, -23, 22, -53, -72, -75, 7, -61, 9, 40, 6, -4, -87, 51, 23, 15, 15, 176, 8, 0, -156, -137, -52, 17, -77, -79, -20, -59, -105, -38, -226, -10, -51, 97, -33, -51, -146, -67, 16, -46, -63, -141, -9, 15, -39, 98, -185, 58, -29, 51, -73, 86, -70, -31, 93, -31, 14, -17, 60, -175, 3, -54, -101, -18, -54, 67, -87, -102, -25, 17, 7, -168, 67, -62, -260, -46, -40, -105, 78, -13, 18, 38, -23, -101, 59, 46, -59, -93, 62, -193, -118, 72, -27, 16, -36, 189, 68, -73, 92, -12, 94, 22, -123, 19, 138, -86, 21, 28, -168, -65, -87, -106, -65, 7, -91, 8, 38, 95, 58, 44, -3, 90, -146, 64, -53, 62, 23, 86, -28, -74, -27, 111, -21, 9, -93, 2, -123, 117, 36, -64, 75, 90, 47, 66, 34, 0, 111, 2, -238, -56, 91, -79, -115, 193, 85, 29, 25, 124, 50, 15, -9, 52, -82, 73, -23, -51, 28, 92, 89, 53, -10, 14, 86, 135, -15, 159, -51, -71, 87, -31, 16, -45, -20, -47, -7, -119, -86, -7, -53, -152, -63, 28, 4, 82, -40, 73, -30, -106, 9, -21, 81, -138, 21, 124, 34, -98, 47, -37, 0, 74, -98, 26, 87, 1, -95, -17, -16, 85, -91, 67, 1, 51, -120, 34, 14, -164, -148, -107, -105, 35, -14, 95, -73, -4, -2, -150, 6, 43, 19, 54, 8, 17, 34, -40, 22, -30, 46, -56, 139, 51, 60, 6, -46, 95, -19, -67, 11, -75, 28, 2, -49, 63, 70, 3, -20, 107, -66, 5, 88, 17, 115, -17, -117, -31, 27, -184, -67, -348, -56, -106, 4, -132, 81, 30, -91, 39, 53, 91, -8, -33, -83, -38, 26, -114, -75, 24, 74, -29, 67, 176, -125, -36, 54, -111, -57, 27, 135, 106, 20, 28, 58, -4, 20, 76, -41, -29, 5, 118, -102, 23, -178, 50, -65, -62, -56, 51, -13, 108, 7, -73, 155, -119, -70, 102, -25, 16, -23, 18, -39, -39, -178, 18, -149, 1, 18, 48, 35, -53, -83, 44, 68, 55, -15, -161, 41, 83, -57, -87, -114, -56, -82, 158, 19, 49, -19, -89, -16, 38, 20, 25, -32, -35, 6, 71, -23, -15, -2, -67, -54, -106, -172, -63, 33, -56, -20, -19, 70, -54, 74, -18, -19, 15, -6, 33, -111, 84, -52, -16, 81, 73, 58, 75, -33, 22, 118, 46, 116, -106, -115, -107, 195, -206, 13, 37, -74, -150, 7, -121, 22, -89, 43, -12, -144, -42, 33, 62, -39, -49, -120, -18, -30, 2, 57, -225, -6, 16, 68, 157, 68, 55, 93, 2, -23, -37, -1, 51, -114, -43, 7, -77, 66, -64, -60, -57, 2, 14, 68, 41, -156, -116, -105, -213, -113, 0, -171, 125, 42, -19, 104, -1, -72, -14, 42, -184, -40, -20, -119, -40, 116, -23, -84, 27, 104, -12, -87, 11, -23, -33, 1, -60, 16, 219, -83, -22, -55, -158, -132, -16, -98, -120, -110, -128, 26, 37, 61, 104, -32, 62, 142, -77, 22, 20, 3, 2, 62, -76, -23, 47, 29, -29, -104, 7, 51, -53, 136, 4, -11, 12, 32, 5, 82, -112, -41, -87, 49, -141, -39, 9, -4, -123, 50, 51, -69, 32, 31, 99, 15, 42, -29, 48, -32, 39, -113, -74, -70, -6, 23, 178, -146, -64, 48, -94, -202, 18, 142, 19, -40, -14, -67, -6, 105, 43, 68, -37, 6, 154, 16, 10, -152, 106, -55, -151, -106, -58, -49, 79, -21, 29, 88, -25, -28, 81, 11, -5, -98, -34, 5, 4, -166, -66, -140, -27, -71, -14, 75, 28, -122, 29, 81, -130, 2, -169, 55, -57, 25, -42, -26, -74, -125, 137, -94, -24, -39, -32, 55, -16, -40, 125, 85, 8, 28, 70, 53, -19, -30, -106, 30, -74, -92, -3, -36, -101, 90, -46, 62, 21, -44, -48, 46, 84, -14, 151, -82, 106, 22, -17, 67, -6, 125, 54, -5, 9, 170, 62, -43, -164, -63, 46, 55, -213, -35, 41, -85, -25, -13, 61, 53, -80, -38, 149, -162, -34, 7, 63, 0, 36, 110, 53, 30, 3, 68, -51, -40, 13, 37, 107, 43, 215, 136, -8, 30, -87, -101, 32, 46, -99, 14, 2, 88, 70, -110, 31, 158, 52, 105, -48, -37, 19, -117, -72, 32, -41, -79, 37, 97, 21, -18, 12, -19, -58, 102, 37, 37, 125, -76, -26, 40, 17, -145, -29, 16, 123, -122, -140, 2, -23, -28, 35, 83, 25, 52, -19, -116, -44, -174, 105, -46, 36, -124, -146, 47, -42, -102, -53, -26, -27, -43, -144, -69, 65, 6, -55, 30, 2, 29, -27, -34, -1, 17, 44, 13, -91, 68, -31, -46, 20, 52, -16, -27, -82, -30, -95, 74, 117, -121, -25, 83, -114, 96, 5, -18, -60, -31, 5, 65, 1, 53, 14, 100, 8, -66, -43, 1, 2, 11, 30, -156, -13, 59, 56, 103, 15, 70, -124, -139, -125, -124, -129, -91, -4, 41, 43, 35, 24, 23, 41, -1, -7, -98, -164, 32, -38, -115, -64, 6, 113, -9, 126, 108, 113, -4, 49, 28, -42, 68, -52, -173, 63, -171, -38, 141, -40, 50, -26, 6, -50, 80, -220, -18, 65, -26, -199, 152, 75, 144, -54, 138, 46, -168, 116, 39, 30, 75, -91, -53, 84, 25, 32, 3, -47, 113, -37, 57, -96, 115, -16, 20, 70, 9, 67, 61, 20, 23, -33, -125, 125, 71, 71, -126, -28, 16, -45, 93, -13, -77, -91, -17, 46, 34, 49, 28, -97, 36, 24, 16, -80, 197, 52, 89, 6, 58, 105, -8, 117, -9, 2, -9, 35, 134, 110, 212, 103, 13, 40, -40, 89, 10, 12, -39, -72, -43, -32, -45, 126, 94, -63, -60, -36, 45, -55, -79, -41, 27, -86, -112, -26, -14, -90, -123, 111, -42, 52, -81, 28, 52, -136, -1, 125, -76, 5, -36, 69, 4, -14, 7, 82, 195, -78, 12, -62, 54, -72, 23, 93, -55, 79, 6, 59, 46, -103, -7, 3, -27, 10, 59, 98, -23, -80, 88, -120, -78, 71, -4, 129, 118, -43, -93, 45, -17, 8, 51, 1, 33, 42, 69, 146, -85, -31, -32, 99, 9, 8, 48, 2, -50, -91, -10, -44, 34, 25, -76, 15, 40, -103, 6, 43, -138, 54, -29, -55, -72, -173, -2, 12, -37, 49, -22, 35, 62, -6, 182, -16, -47, -43, -67, -93, 140, -77, 23, 94, 110, 11, 97, -1, 200, 51, 21, -11, -24, -114, -40, 198, 126, 96, 183, 65, 66, 76, -120, -97, 7, 62, -109, 21, -30, 14, 75, 37, 62, 157, 31, 149, 14, -99, 18, -85, -25, -56, -10, -46, 23, 83, 71, -39, 105, -47, 56, 0, -2, 2, 35, -2, -19, 70, 13, 31, 62, -36, 92, 28, -133, -17, -74, 18, 64, 4, 81, 19, -70, -63, 4, 79, 116, -89, -3, -29, -71, 90, -57, -33, -62, 109, -131, 46, -72, -92, 91, 8, -73, 51, -57, 6, 70, -106, 6, -2, 47, -32, 19, -15, -30, -60, 29, 198, -50, -48, -45, 15, -180, 51, -262, -28, 32, 45, -97, 70, 83, -14, -16, 9, 78, 152, 60, -61, -51, -13, 87, -34, 45, 15, -47, 96, 223, -47, -45, 82, -83, -90, -27, 169, 18, 36, -46, 25, -26, -14, 99, 40, -20, 37, 91, -31, -34, -124, 93, -60, -146, 6, -71, -4, 46, 1, 98, 25, -14, 148, 22, -20, 8, -69, 21, -75, -78, -100, 85, -157, 93, 23, 59, 15, -35, -9, -38, 201, -33, 39, -100, 40, -55, -11, -109, -85, -97, -133, 150, -74, -24, -115, -50, 67, 65, 114, 187, 71, -89, 41, -24, -83, 22, -30, -82, 34, -17, -62, -79, -27, 28, 184, 41, 96, -73, -38, -52, -19, 77, -64, 68, -128, 6, 49, 4, 9, -12, 106, -32, 57, 76, 128, 7, 147, -164, -62, -31, -131, 68, -39, -9, -34, -7, 12, -81, 36, 26, 4, 78, -48, -100, 2, 22, 42, 46, -71, -76, 47, 95, 203, 67, 26, -28, 48, -112, 24, -68, -47, 25, -60, -93, -29, 35, -52, -93, 20, -11, -47, 22, 78, -3, 26, -63, 55, -39, -176, 14, -122, -199, 132, -68, -36, 103, -39, 119, -16, -93, -124, -33, -21, 36, -42, 60, -123, -93, 72, 12, -48, -38, 159, 21, -74, -45, -14, 43, 41, 61, -8, 76, 61, 70, 69, -42, -139, -61, -37, 6, -92, -124, -8, -19, -37, -25, 66, -30, -5, -120, 10, 27, -46, -70, 52, -6, 81, -83, 55, 89, 38, 49, -8, 4, 64, 69, -14, 73, 161, -6, 5, -43, -44, 14, -61, -226, -67, 29, 124, -180, -22, -94, 9, 115, -15, 32, -1, 29, -16, 44, 116, 115, -25, -41, -88, 7, 1, 5, 34, 5, 4, 19, 153, 34, 49, -81, -100, -112, 41, -60, -10, -19, 106, 19, 35, 95, 25, 157, 56, -24, 23, 73, 5, 26, 11, -14, -48, 95, 188, 48, 137, 108, -38, 169, -132, -19, 10, -14, 48, 43, 21, -2, 175, 21, -26, 134, -56, -138, -8, 69, -7, -82, 122, 51, -72, 141, 29, -70, 17, 59, -178, 38, 40, -2, 63, 85, -63, 104, 189, 130, 133, -85, -14, -32, -101, -43, -130, -65, -18, 6, -6, 7, 98, 12, 33, -2, -38, -1, 19, 36, -35, -41, -84, -41, 12, -31, 27, -24, -35, 14, 80, -73, 165, 17, 382, -68, -132, -129, 117, -67, -74, 37, 78, -26, 57, -127, -66, -33, 87, -92, -43, -65, 135, 15, -65, 46, -58, -10, -11, -17, 58, -226, 57, -7, 105, 125, 50, -42, 13, 78, -10, 49, 38, 95, -143, -37, -45, -83, 53, -21, 62, -103, -63, 90, -20, 61, -167, 26, -102, -159, -49, -40, -121, 76, 29, 32, 64, 15, 4, -24, 10, -52, -5, -17, -101, -66, 30, 5, 151, -6, 133, 48, 119, 79, -133, 15, -34, -84, -19, 109, -10, -32, 39, -132, -86, -72, -7, -124, -73, -118, -2, 22, 70, 79, 46, 44, 93, -112, -17, -11, -41, 6, 91, 4, 16, -3, 81, 7, -33, -27, 22, -68, 98, 7, 35, 22, 93, 36, 11, -8, 3, 74, 51, 18, -33, -11, -30, 219, 0, 30, -2, 30, -103, -15, 137, -26, -2, -37, -18, 43, 162, 162, 31, -2, 13, -18, -46, 42, -15, -57, -1, 33, -28, -32, 175, -6, 79, -11, -113, -17, 82, 63, -9, 30, 40, -58, 78, -34, -128, -128, 150, -10, 152, -134, -19, 78, -112, 83, 138, -109, 58, -65, -24, -128, -67, 48, -39, 124, -90, 3, -31, 111, -79, 0, 149, -94, 50, -47, 12, 6, -78, -66, 75, -3, 32, -9, 46, 10, -71, 35, -25, -58, 95, -109, 43, 58, -46, -132, -27, -23, 7, -26, 56, -150, 118, -32, 115, -30, -34, 4, 77, -45, 96, -1, 30, 36, -59, 10, -55, 24, 35, -104, -38, 83, -135, -111, 52, -56, 61, -35, 15, 4, -48, 109, 87, -22, -53, 156, -25, 42, 165, 25, -21, -18, 19, 63, 70, -113, 174, -11, 103, -32, 87, -35, -25, 85, -58, 37, -147, -44, 30, -96, -85, -1, -11, -187, -81, 37, -42, -5, -50, -110, 22, 49, -123, -46, -51, -20, 44, -50, -107, 13, -121, 29, 76, -24, 29, 99, -34, 6, 49, -101, -141, -71, -49, 92, 84, 145, -125, -41, 21, -73, 68, -5, -43, -28, 96, -38, -89, -106, 29, 0, 5, 10, 10, 1, -46, -134, -89, -59, 26, 110, 120, -32, 125, 18, 139, 129, 2, 55, 83, -15, 39, 44, 33, 83, -4, -64, 19, 58, -82, 55, 3, 15, -7, -24, 20, 15, 48, -10, -48, -8, -2, -1, -104, 19, -96, 130, -24, 4, -37, 105, 55, -62, -105, 21, 195, 9, -61, 70, 62, 62, -78, -104, 61, -9, -119, -58, 10, 46, 94, -71, -10, -25, 64, 119, -21, 37, 130, 68, -40, 24, -69, 95, -244, -96, -25, 18, -52, 76, 29, -83, -21, -90, -25, -77, 3, 71, 2, -199, -22, -50, 91, -64, -35, -30, 0, -41, 21, -21, 60, 59, 39, -1, 20, -32, 52, -85, -63, 7, -63, -67, 90, 10, 5, 139, 7, 85, -111, 105, 125, -109, 82, 39, -60, -73, 43, -93, -12, 76, -133, -9, 10, -35, -143, 57, -28, 50, -42, 79, 50, 22, 23, 13, -59, -7, 32, -100, 10, 63, -15, 66, 74, -21, 17, -124, 6, -71, 83, -32, -59, 48, -9, 60, 14, 10, -8, 41, -77, -95, -393, -111, -124, -64, 104, -118, 6, 28, 130, 40, 42, -40, 0, -129, 0, 33, -139, 71, 236, 5, -11, 33, -24, -1, -49, -52, -6, -280, -26, -6, 82, 199, 38, 135, 5, 80, 41, -101, -133, 7, 55, -112, 59, -66, 44, 69, -31, 9, 73, 123, 62, -34, -65, 30, -152, -65, -95, 7, -43, -39, 44, -38, 78, 30, -11, 48, 74, -129, 3, 31, 30, 21, 129, -13, 175, 3, -83, 85, 134, -126, -44, -113, 20, -24, -18, 141, 60, -57, -151, -51, -203, 33, -5, -86, -166, -56, 87, -24, -3, 1, -17, -95, 36, -108, -53, -36, -152, 0, 53, -1, 42, 8, 1, -65, -26, 25, 76, -46, 90, -33, -47, 58, -17, -71, 47, -47, -79, 24, 138, 51, 81, 59, 74, 196, -178, 26, 80, -19, 3, -28, 91, 66, -43, -52, 118, 26, 51, 19, 7, -10, -19, -35, 63, -66, -78, -110, -144, -43, -6, -65, 146, -59, 231, 152, 23, -1, -57, -30, -38, 87, 27, 69, 125, -17, 71, -49, 84, 212, 86, 62, 41, -39, -83, 0, 71, -3, 62, -56, 6, 0, 42, 50, 65, 8, 110, 8, 45, 0, -71, 155, 65, 50, -44, -63, 68, -114, 72, -92, -113, 150, -105, 70, 131, -47, 1, 63, -21, -50, 80, 37, 36, -111, 47, -91, -41, 10, -32, -77, -16, -21, -48, 37, 66, -23, -16, 69, -105, -83, -26, -23, -15, -84, -38, 45, 39, -31, 62, 0, -41, 5, -19, -56, -99, 6, -75, -58, -65, 84, 161, 141, 48, -120, 34, 124, 60, 54, 172, 170, 26, 42, -65, -41, 2, -92, 157, 6, 155, -14, 7, 48, 77, 24, 2, 33, -70, -149, -44, -87, 43, 119, 26, -46, -22, 101, 7, -113, -59, -110, 151, 7, -81, -58, -13, 43, 60, 21, 20, 25, -14, 37, -5, -63, -67, 49, -40, 129, -11, -72, 20, -39, 8, 50, 76, 7, -48, -68, 9, -64, 87, 74, 92, 99, 89, 57, -122, -99, 97, -120, -80, -141, 38, -10, -90, 49, -67, -106, 4, 88, -33, 97, -22, -18, -52, 103, 102, -6, 96, -71, 34, -32, 61, 102, -41, 19, -126, -65, -6, -51, 23, 85, -52, -3, -57, 150, 51, 67, -21, -112, -8, 68, 14, -1, -32, 90, 56, -55, 103, 53, -170, -90, 40, -252, 221, -33, -68, 54, 16, 83, 64, -7, 21, 2, 125, -33, -57, 13, 37, 96, 114, 60, -141, -20, 119, 19, 104, 44, 8, 66, -93, -85, -91, -61, 38, -3, 7, -80, 18, 83, -107, 74, -17, 83, 5, -30, -76, -108, -83, 6, -58, 53, 119, 37, 33, 155, -87, 54, 5, -51, 66, -71, -206, -31, -166, -54, 144, -41, 112, 21, -110, -6, 66, -23, -34, -45, -39, 61, -23, -33, -12, -95, 73, 85, -80, 67, -74, -42, 73, -112, -24, 154, 79, 5, 116, -37, 51, 9, -69, 35, -78, -100, -154, 15, 44, -87, 117, 19, 90, -1, -52, 22, 102, 135, -54, 26, -78, 76, 85, 12, 95, 45, 13, 100, 103, -11, 200, -41, 121, 60, -7, 67, -25, 42, 29, 25, -16, -125, -27, 19, 56, 37, 61, -174, 124, 56, -101, -102, 37, -119, -64, -48, -6, -63, -58, 84, 77, 48, -171, -127, -96, -156, -98, 14, -82, 91, 90, -29, -89, 124, -68, 50, 1, -67, -68, -25, -139, -54, -107, 41, 131, 25, 60, 103, -16, 42, 76, -70, -115, -120, -8, -82, -28, 20, -27, -2, -15, -65, -15, -17, -36, -12, -146, -23, -18, -79, -68, 114, 51, 83, 16, -56, -10, -87, -129, 51, 77, 36, 141, -63, 71, 28, 102, 69, -60, 64, 79, 53, -64, 87, -21, 125, 81, -114, 108, 75, -67, 37, -103, -33, 0, 36, 39, -54, -34, 7, -76, 82, 36, -72, -215, 63, 0, 24, 34, 138, -19, -112, 32, 64, 35, 51, 9, 185, 37, -39, 9, 11, 158, 49, -49, -77, -35, 87, 22, -57, 81, 4, -7, 26, 73, -8, 53, -197, -151, -52, 5, -26, 29, 35, -22, 14, -34, -24, -11, -91, -90, 22, -27, -95, -122, 11, -3, -152, -9, -138, -55, -16, 33, 160, -206, 36, 135, -104, -62, -78, 15, -15, -61, -8, 108, 172, -33, 22, -122, 23, -20, -73, 30, 39, 110, -234, 114, -64, -138, -176, -14, -62, -100, -23, -45, -16, 26, -105, -81, -41, 93, 107, 159, 99, 27, 64, -22, 88, 15, 72, 34, 3, 107, 123, 71, -49, -39, 38, 38, -28, -17, -78, 9, -81, -28, -78, -7, 84, 81, -21, -7, -31, -3, -94, 91, -117, 69, 92, -181, -11, -275, 5, 7, -79, -66, 150, 4, 70, 137, 7, -65, -156, -100, -43, 72, -44, 170, -112, 11, 18, 97, 3, -92, 71, -28, 49, -2, -179, 39, -153, 15, -47, 63, -116, -52, 114, -33, -21, -133, -118, -122, -63, -37, -1, -62, 59, 198, -88, -24, -39, 13, -11, -75, 81, -114, -98, -23, -40, -26, -14, -48, 28, 46, 139, 3, 194, -52, -8, -51, -27, 26, 33, 102, -36, 183, 19, 46, -83, 88, -128, -87, -9, 80, 26, -82, -5, -24, -52, 112, -53, -28, -77, -18, -30, 20, 81, -43, 11, 80, -93, 198, -58, 63, 44, -28, 26, -17, -43, 13, -25, 72, -21, -70, 53, 16, 93, 30, -42, 31, -92, 2, 92, 160, 19, -26, 90, -55, 33, 65, 257, 69, 49, 82, -108, 52, 2, 57, -88, 26, -6, 6, 69, 33, 34, -88, -25, -60, -200, -95, 54, -95, 88, -168, -33, -31, 52, 42, 81, -18, -119, -153, -90, -67, -108, 25, -81, -15, 7, -38, 97, 152, 3, 39, -73, 17, -21, -61, 73, -147, -72, 41, 106, -20, 78, 23, -7, 119, 27, -48, -215, -54, 31, -141, -60, -30, -85, 25, -36, -35, 71, -11, -41, -24, -227, -53, -90, -21, -141, 156, 70, -6, -20, 27, -14, -47, -68, 97, 62, 128, -35, -147, -15, 46, 35, 30, -44, 132, -56, 2, -31, 38, -73, 146, 121, -8, 1, -85, -116, 7, 40, -45, 40, 11, 9, -1, 65, 85, -34, -11, -37, 35, -120, -77, 67, -37, 71, 116, 24, -68, 69, 20, -16, 160, -214, 12, 5, -88, -58, -63, -84, 54, -44, -69, 20, -56, 47, -89, -17, -48, -102, -17, 120, 16, -82, 7, 108, 22, 26, -19, 16, 50, 193, 136, -65, -24, 0, 79, 80, -38, 62, 71, 132, -67, 72, 41, -22, 175, 8, 81, -4, -26, -29, 17, -95, -48, -7, -21, -15, 78, -6, 29, 169, -85, 170, 10, -34, 31, -51, -34, 62, 11, -104, -49, 49, -19, 116, -101, -73, 140, -86, 41, -68, -106, 95, -53, 72, 28, -43, 46, -62, -172, -10, 60, -122, 17, -23, 8, -12, -16, -77, 27, -42, 24, 45, 30, -77, 1, -96, -4, 80, -78, -9, -61, 41, -90, 94, -9, -119, -51, 20, -91, -89, -22, -102, -1, -92, 50, 86, -37, -63, 45, -78, -16, -88, 5, 37, -9, -21, -17, 45, 5, -1, 17, -1, -9, 86, -81, 29, -22, 78, -190, -26, 6, 55, -63, 17, 8, 2, -75, -53, 6, -90, -10, -53, 45, 53, 47, 113, 93, 83, 39, -13, -67, 74, -108, 109, 23, -108, 2, -70, 145, 51, -79, 41, 116, 1, -1, -59, 17, 5, -211, 13, -84, -89, 122, 7, -43, 154, -66, -72, -24, 153, -100, -63, 110, 201, 110, 89, 50, -20, 93, 80, -24, 29, 47, 2, 85, -164, -160, -13, 49, -131, 29, -75, 96, -20, 64, 12, -26, -133, -44, 32, -26, -118, 10, 1, 86, 81, -77, 60, -54, 24, -21, 19, -13, 7, 25, -42, 22, -71, -48, 31, 9, -18, 236, 46, -295, 69, 165, 38, -173, 121, -51, -42, 60, 94, 15, 51, -100, 99, -51, -13, 66, 93, -27, 38, 15, -58, 23, 162, 53, 2, -96, 299, -16, 12, -42, -132, -47, -26, 29, -53, 23, 51, 91, -57, 9, 40, 84, 68, 2, 24, 134, 127, -18, -45, -53, -29, 108, 143, 61, 153, 65, -73, 166, -77, 45, 11, -96, 185, 33, 67, -82, 87, -9, -33, 21, 40, -116, -54, 150, 40, 18, -9, 123, -104, 45, -13, 26, -56, -7, -142, 30, -22, 69, 6, 152, 27, 75, 78, 219, 87, 10, -61, -77, -102, 30, -68, -30, 37, 13, -7, 114, 58, 30, 11, -58, -26, -10, 29, 14, -55, -89, -43, -71, -79, -27, 30, -7, -47, -11, 55, -17, 89, -1, 316, 45, 23, 25, 88, -109, -83, 38, 97, -99, -57, -16, -76, 45, 62, 6, 164, 157, 83, -42, 2, -11, -131, 115, -55, -49, 92, -54, 38, -42, -104, 1, 44, 40, -24, 11, -46, 55, 75, -6, -54, 19, 19, 180, -51, -28, 82, 73, 3, 111, -69, 20, 59, 103, 81, 23, -44, -32, 49, 43, 19, -67, 49, 188, 76, 155, -19, 60, 15, -76, 49, 83, -46, -126, 173, -68, 129, 138, 138, -34, 102, 50, 88, -25, -42, -15, 41, 21, 10, -17, 36, -31, 57, -5, 70, 126, -56, -36, 42, -44, 85, -15, 15, 55, 4, -85, 66, 71, 57, 43, -40, -53, 86, -50, 30, -75, -57, -87, -79, -19, 35, -19, -46, -5, -20, 111, -64, 79, 53, -27, 126, 31, 2, 132, -17, 107, -33, -117, 79, 7, -40, -33, -49, -34, -169, -79, -9, -68, 36, -3, -67, -10, 87, 20, -72, -64, -62, 21, -18, 90, -14, 55, -1, 55, 10, -49, -73, 15, 34, -16, 35, -80, -5, 13, 80, 21, -31, -43, -97, 69, 36, -54, -126, -83, -40, -167, 5, -61, 32, 82, 12, 28, 108, -59, 24, 45, -247, -63, -61, -132, 39, 122, -79, -36, 116, 28, -161, -103, -4, -96, -94, 61, -189, -40, 153, -115, 65, 83, -114, 75, 1, -124, -124, 37, -108, 104, 6, 51, 48, -37, -27, 124, -46, 43, -5, 42, -76, -46, -105, -70, 107, -127, 59, -156, 47, -45, 100, 12, 29, -1, 73, -6, -55, 22, -127, -5, -148, 11, 130, 122, 22, 88, -71, 149, 16, -104, 22, 57, 9, 85, 42, 103, 4, -52, 89, 94, -98, -43, -71, 40, 128, 5, 53, -49, -120, 265, 14, 97, -98, -112, -100, -83, -47, -98, 52, 106, 117, 70, 81, 18, 0, 70, -33, -57, -58, 87, -60, -9, -94, -11, 96, 43, 168, 202, 108, 8, 105, -78, -62, -4, -83, -69, 2, -105, -26, 148, 55, -35, 38, 0, -112, 7, 8, 27, -96, -52, 46, 107, 37, 62, 7, -20, 52, -118, 29, 34, 28, 92, 204, 24, 85, 85, 103, 39, -17, -30, -51, 54, -77, 72, -118, 97, 56, -50, 124, -17, 24, -7, -48, -51, 36, -12, 15, -65, -59, 72, -130, 0, 57, -52, -123, 42, 14, -23, 24, 98, -69, 164, 102, 48, -66, 85, -10, -51, 19, 133, 103, -58, -138, -97, 49, 57, 47, 45, 96, 112, -7, -5, -24, -61, 86, -13, -38, 135, 70, -1, -92, -22, 31, 0, 3, 38, 47, -34, -72, 67, -19, 44, 37, 97, 199, -104, 75, 158, 73, 64, 63, -66, 16, -77, 148, -16, -16, 35, 92, 103, -57, 40, 51, 51, 215, 21, 122, -53, 71, 2, -79, 115, 36, -67, -143, 258, -38, -32, 72, 223, -50, 93, -30, 113, 82, -114, 2, 85, -6, 40, -15, 12, -66, -31, -62, 35, 70, -33, 6, 28, -8, 91, -79, 22, 83, -22, -43, -63, -51, 8, 2, 29, -2, 20, -76, -60, 41, -32, 50, -82, -106, -37, 17, 10, -49, 40, 75, -110, 98, 60, 209, 37, -9, 8, -123, 138, 34, -25, -21, 26, -15, 2, 31, -8, 70, -91, -39, -61, -176, -49, 54, -90, 102, -173, -15, 56, -25, 23, 6, -29, -5, -147, -92, -81, -104, 14, -29, -39, -24, -10, 80, 119, -46, -54, -50, 41, -98, -80, 11, -173, 0, 69, 57, -17, 11, -22, 40, 135, -35, -51, -211, -72, 29, -173, -103, -53, -109, -19, -18, 3, 110, -53, -26, 0, -252, -35, -194, -63, -110, 131, 12, 17, 30, 35, 52, -33, -47, 92, 92, 26, 29, -179, -69, 59, -17, 58, 15, 88, -39, -16, -29, 86, -98, 80, 69, -4, -19, -116, -128, -47, 53, -53, 29, 77, 3, 8, 56, 96, -11, 28, -42, 37, -115, 24, 74, -26, 93, 67, 22, 89, 27, -58, -84, -80, 84, -109, -1, 115, 21, -52, -217, -32, -70, 49, -39, 48, -113, 38, -3, 71, -7, -125, 79, -55, -25, 76, -154, 49, -116, 91, 16, 69, -39, 1, 160, 8, -91, -77, -68, -145, -63, -20, -11, 24, 98, 232, -85, 56, 22, 31, -39, -146, 118, -84, -193, 31, -88, 36, 4, 27, 26, 28, 157, -31, 184, -72, 7, -114, 61, 13, -60, 129, -95, 219, -69, -20, 15, 128, -118, -71, -73, 47, -28, -144, 89, -55, 54, 81, -110, 27, -157, -102, -19, 99, 50, -49, 12, 38, -103, 220, -108, 15, -71, 67, 37, -72, -101, 5, -71, 38, 34, -41, 63, 84, 55, 3, 5, 116, -27, -84, 137, 177, 32, 3, 73, -40, 42, 65, 85, 177, 108, 52, 191, -176, 93, -15, -78, -5, -14, 116, 17, 38, -79, 3, -85, 133, -82, -16, -32, -14, -8, 151, 30, -91, -77, 207, -46, 27, -70, 95, 4, 111, 79, -105, 22, 4, 82, 53, 12, 61, 49, 162, 25, 50, -55, 161, 78, 15, 25, 31, 110, -147, 34, 162, -67, 47, 61, 31, 40, -84, 28, 168, 53, 82, 12, -53, 29, -48, -35, 174, -71, -102, -57, 62, 34, -64, -87, 20, 59, -25, 26, 38, -76, -27, -81, 69, 31, 53, 87, 138, -54, -9, 87, -138, 22, -41, -1, 45, -97, 13, 44, 35, -72, -33, 119, -2, -38, -36, -102, 66, -64, -59, -122, -10, -58, 77, -47, 2, -9, -83, -59, -17, -35, -114, -4, -186, -66, 32, 126, -2, -58, -51, 65, 3, 36, 32, 49, -63, -198, 2, -39, -43, -55, -14, -133, 1, 27, 64, -67, -126, 48, 26, 44, 94, -31, 0, -181, 69, -46, 39, -61, -17, 86, -84, -80, -42, -106, -44, 11, -97, 89, -100, 111, 96, -26, -2, -81, 47, 40, -24, -64, -101, -97, -22, 40, -30, 55, -35, 80, 85, 153, -69, 81, -134, -71, -90, 17, -38, 39, 80, -119, -24, 22, -7, -131, -75, -38, -38, -33, 55, 61, -183, 85, -46, -7, 115, -38, -24, -86, -179, -72, 106, -88, 23, 36, 54, -1, 155, 33, 92, 82, 50, 14, -37, -148, -15, -131, 74, 51, -47, 76, -66, 73, -52, 118, 32, -31, 14, 54, 105, -94, -32, -44, 17, -145, -32, 527, 44, 33, -117, 248, -6, 82, 120, -30, -54, -8, -4, 75, 38, 39, -141, 174, 21, -4, 61, -29, -71, -103, 79, 28, 6, -13, -210, 77, -101, -32, 106, 113, -3, 21, 8, -42, 20, 27, -14, -94, 25, -129, -90, 15, -12, -142, -9, -110, -22, -58, 61, 29, -237, -48, 30, -145, 67, -119, 51, -121, -10, 92, 156, 98, -20, -22, -163, -77, -81, -60, 119, 82, 93, -158, 25, 62, -144, -186, 71, -117, 11, 51, -39, 12, 84, -121, -61, 55, -34, 61, 55, -13, -76, -38, 10, 6, -30, 169, 97, -14, 125, 179, 158, 41, -91, -7, -24, -14, -40, -82, 68, -47, -18, -39, 11, 56, 124, -61, 11, 70, -44, -109, 71, -80, 77, 81, -154, -3, -23, 0, 86, 129, -169, 33, 29, -47, -66, -40, 18, 160, 57, 29, 35, 126, 125, -13, -78, -62, 88, -7, 24, -46, -31, 28, -121, 80, -8, -10, -114, -73, -96, -40, -37, -42, 36, 36, -102, -46, -7, -35, 87, 12, 25, -73, -123, 58, -36, -94, -42, -104, 148, -96, 107, 150, 41, -51, 31, -65, -37, 11, -53, -4, 95, -24, -8, 130, 16, 51, 41, 30, -127, 37, -188, 1, -26, 12, -154, -65, 110, 69, -25, 163, -25, -238, 75, -80, -91, 160, -8, 72, 120, 128, 60, 124, -43, 14, 31, -76, -41, -7, -44, 71, 23, -20, 49, 64, -11, 27, -20, -86, 8, 34, 137, -101, 1, -90, -13, 38, 6, -79, -99, 51, -72, 36, 51, 46, 14, -410, 17, -7, -10, 2, 52, 21, 7, 2, -66, -35, -81, -77, -108, -156, -42, -59, -47, -49, -63, -54, -44, -16, 18, 26, 12, -18, -1, 17, -4, 12, 16, -37, -22, -47, -67, -127, -130, -162, -156, -174, -167, -264, -198, -147, -109, -127, -167, -132, -151, -125, -103, -74, -6, 11, -11, -3, -7, 7, 3, -28, 16, -14, -3, -40, -85, -87, -109, -117, -96, -88, -90, -107, -68, -77, -59, -138, -89, -81, -64, -53, -22, -17, 16, -17, 15, 31, 17, -11, -35, 1, 31, 14, 14, -9, -60, -73, -73, -41, -58, -56, -70, -3, 0, -26, -45, -13, 19, -39, 5, 1, -16, 15, -1, 69, 21, -52, -100, -57, -8, -10, -28, -46, -72, -53, -30, -27, -28, -27, -35, -6, 24, -18, 16, 14, 29, -29, -40, 47, -14, -8, 7, 61, -17, -79, -133, -70, -36, -61, -32, -31, -24, -10, 4, -11, 8, -13, -17, 2, -13, -25, -28, -13, 2, -42, -78, -28, 23, 7, -2, 24, -84, -118, -107, -102, -102, -95, -43, 13, 37, 7, 22, 31, 27, 23, 0, 26, 7, -19, -6, -30, -21, -90, -35, -24, 0, 24, -8, 5, -77, -134, -125, -140, -123, -69, -74, 7, 33, 31, 40, 72, 55, 42, 40, 49, 46, -18, -21, -46, -42, -41, 3, 15, -16, 10, 21, 2, -39, -65, -101, -89, -69, -89, -72, 3, 14, 24, 21, 38, 57, 75, 62, 21, 16, -16, -13, -35, -51, -54, 34, 34, -3, 6, 0, -36, 8, -12, -77, -94, -34, -87, -42, -21, -16, 12, 20, 45, 59, 40, -18, -36, 9, -10, -55, -50, -54, -31, -3, -52, 9, -35, -13, -56, 1, -36, -47, -32, -42, -34, -27, 14, -20, -22, 7, 35, 23, -12, -37, -24, -25, -10, -11, -9, -13, -17, 6, -15, 38, -17, -3, -74, 29, 10, -9, -14, -5, 2, 9, -10, -17, -9, -3, 38, 56, 0, 5, -33, -15, -27, 2, 42, -5, -30, 26, 16, 5, -28, -5, -91, 20, 26, 27, 50, 53, 46, 54, 19, -6, 3, 27, 39, 18, 6, 5, -12, -5, 17, 35, 63, 40, -41, 0, 30, 13, 17, -32, -86, -9, 52, 45, 76, 50, 89, 57, 23, 15, 33, 28, 11, 10, 17, 19, 41, 58, 61, 65, 82, 94, -23, 41, 17, 1, 31, -27, -72, -11, 78, 73, 59, 70, 48, 22, 25, 13, 51, 34, 11, -8, 23, 46, 60, 58, 56, 73, 86, 84, -19, 35, 13, -33, 16, 2, -18, -24, 25, 67, 54, 41, 44, 11, 17, -17, 47, 51, 41, 81, 65, 36, 52, 37, 55, 48, 51, 18, -59, 48, -14, -21, 4, 1, -43, -51, -12, 41, 48, 40, 18, 34, 27, -4, 67, 81, 67, 49, 19, -24, -14, 2, -25, 3, 7, -2, -42, -23, -19, 32, -5, -31, 3, 20, 46, 10, 13, 5, 19, 28, -4, 45, 56, 104, 9, 11, -35, -62, -44, -43, -26, -20, -61, -44, -40, -17, -22, 24, -13, 17, -17, 2, 45, 13, 7, 0, 9, -43, -48, -12, 8, 22, -22, -68, -85, -69, -122, -95, -23, -31, -66, -38, 48, -23, -32, -2, 0, -48, -60, 9, 8, -3, -30, -43, -32, -59, -84, -35, -71, -81, -89, -80, -90, -94, -90, -43, -64, -29, -40, 6, 52, 3, -24, -18, 16, 16, -14, -10, 28, -11, -30, -106, -120, -109, -98, -88, -82, -63, -44, -78, -83, -69, -74, -69, -33, -6, -45, 54, 61, -33, -43, 21, 15, 8, -15, 3, 53, 32, -51, -81, -84, -101, -76, -84, -48, -50, -29, -53, -64, -82, -98, -44, -56, -47, -20, 11, 33, -22, -32, 28, 19, 39, -7, -11, 53, 43, -19, -17, -41, -58, -83, -77, -32, -17, -27, -31, -64, -50, -35, -52, -16, -19, -16, -20, 43, -16, 23, -11, -2, 34, -14, -57, -63, -4, 3, 32, 8, 18, -4, -66, -87, -43, -33, 10, -22, -71, -42, -43, -33, -18, -24, 28, 21, -35, -12, 14, -4, -20, -19, -46, -16, 7, -16, -37, 3, 28, 34, -17, -17, -5, -32, 9, -46, -3, 3, -3, 14, 35, 32, 32, 8, 0, -10, 4, 7, 4, 5, 5, -14, 58, 12, 36, 39, 38, 17, 9, 23, 35, 48, 21, 48, 29, 4, 14, 20, 45, 44, 21, 25, 10, -3, 17, 6, -7, 1, 17, 4, 29, 74, 49, 37, 31, 42, 16, 14, 26, -18, 3, 61, 27, 27, 38, 38, 61, 57, 9, 13, -4, 13, -6, -16, 1, 18, -17, 0, -18, 19, 3, -10, 17, 13, 19, -19, -12, -15, 32, 6, 5, 1, -4, 18, 0, 6, -17, 4, 6, 11, 12, -12, -1849, 0, 6, 13, 0, 25, -25, -46, -33, -18, -21, 11, 43, -7, -52, 9, 7, 5, 26, 15, -19, 3, 8, 25, 9, 11, 20, 1, 17, -20, 8, 18, -25, -55, -36, -64, -68, -34, -62, -76, -37, 18, -12, -40, -68, -18, -23, -2, 18, -31, -77, -85, -91, -4, -19, 2, 4, -9, 37, 21, -28, -50, -118, -112, -102, -124, -119, -55, -6, -11, -15, -4, 3, 5, -44, -22, -39, -50, -77, -40, -19, 34, -30, 5, -18, -16, 34, 38, 42, -49, -72, -66, -77, -81, -75, -17, -15, -22, -5, 9, -25, -16, -45, -39, -28, -22, -12, 12, 17, 11, 3, 9, 2, -15, 62, -5, -9, -25, -29, -23, -34, -11, -45, -55, -18, -22, -54, -15, -31, -16, 15, 18, -7, -1, 13, 55, 60, -16, 27, 7, -18, -14, 48, 25, 1, -26, 6, 1, -31, -19, -28, -24, -9, -18, -15, -29, 14, 1, 29, 53, 50, 19, -5, 29, 24, 23, 34, 14, 18, 7, 40, 53, 13, 29, -25, -15, -6, -4, -14, -28, -17, 14, 34, 39, 10, 11, 28, 45, 49, 37, 31, 43, 12, 11, 31, 8, 17, 3, 43, 21, -24, 0, -7, -7, -39, -69, -57, -12, 25, 31, 80, 26, -4, 25, 22, 55, 33, 72, 60, 39, 89, 43, 36, -25, -15, 38, 37, 94, -2, -16, 6, -28, -34, -41, -24, 22, 51, 83, 59, 47, 38, 36, 36, 22, 31, 47, 40, 31, 70, 39, -4, -17, -16, 40, 84, 107, 38, 14, -8, -21, -52, -25, 18, 58, 74, 41, 44, 42, 77, 5, 21, 4, 24, 62, 13, 20, 63, 64, 14, 2, 34, 41, 35, 100, 5, 10, -5, -21, -38, -21, -3, 20, 12, 27, -4, -1, 26, 9, -6, -16, -9, -3, 30, 16, 7, 56, -5, 0, -15, 64, 50, 59, 25, 14, 1, -6, 17, 24, 1, 13, 27, 20, 16, 66, 37, 13, -3, 2, 6, -7, 31, 35, 14, 27, 10, -11, 7, 18, 41, 42, 55, 15, -24, -6, -3, 19, 9, -13, -14, 11, 36, 66, 43, 17, -1, -30, -9, -17, 16, -25, -74, -32, -44, -6, 12, 46, 39, 36, 10, 40, 5, -16, 3, 27, 20, -7, 28, 18, 49, 53, 31, 15, -24, -58, -60, -56, -55, -66, -147, -54, -9, -31, -3, 18, 31, 49, 60, 44, -32, -15, -8, 0, 24, -1, 12, 9, 9, 16, -41, -79, -125, -125, -115, -153, -129, -128, -129, -64, 34, -16, -5, 25, 17, 4, 6, -31, -32, 13, -5, -14, 11, -26, -15, 13, -5, -70, -128, -168, -189, -197, -117, -119, -141, -119, -87, -75, -12, -24, 25, -23, -60, -43, 7, 18, 8, 55, -9, 6, 5, -4, 19, 6, -4, -100, -175, -192, -146, -109, -41, -37, -81, -32, -72, -55, 1, 18, -4, -7, -11, -2, 5, 37, 22, 36, 42, 27, -1, 26, 18, 42, 1, -98, -159, -104, -25, 10, 47, 17, -6, 20, -10, -41, 33, 44, 8, 7, -38, -62, -38, 7, 10, 28, 22, -4, -6, 15, 8, 74, 31, -50, -71, -41, -1, 35, 26, 24, -9, 35, 69, -10, -1, 55, 27, -22, -55, -78, -87, -22, -23, -14, 12, -17, -20, 4, -27, 22, 20, -46, -25, 29, 39, 53, 31, 9, -36, 41, 58, -26, -9, 50, 29, 3, -24, -80, -61, -52, -32, 11, 18, -26, -33, -38, -28, 0, 13, -31, -3, 17, 27, 27, 42, 22, 1, 10, 71, 14, -5, 46, 8, 14, -31, -61, -29, -80, -53, -48, -25, -27, -32, -35, -1, -39, -35, -57, -12, 3, 46, 8, 1, 21, 13, 49, 73, 24, 2, 27, -5, 21, -38, -61, -6, -27, -41, -53, -13, -16, -27, -45, 14, 6, -26, 1, -46, -6, 21, -12, 18, -16, -2, 56, 46, 4, 22, 4, -19, 10, -29, -22, -29, -31, -24, -52, -39, -12, -2, -39, -39, 3, 10, 5, -48, -22, -39, -25, 17, 12, 41, 34, -5, -37, 1, 10, -7, -9, 29, 12, 43, -3, -36, 15, -16, 23, 2, 30, 56, 40, 48, 33, 55, 54, 7, 62, 68, 73, 36, 26, 10, 34, 9, -2, 20, 10, 11, 64, 80, 84, 44, 93, 44, 48, 45, 62, 74, 91, 52, 44, 118, 124, 94, 133, 108, 52, 47, 16, 52, 0, -12, -11, 3, -13, 6, -8, 0, 32, 49, 42, 77, 64, 110, 70, 65, 58, 12, 32, 54, 38, 38, 33, 58, 56, 27, 22, 15, -2, 7, 4, -15, 0, -17, -20, -12, -14, -10, -9, -19, 0, 6, 4, 21, -4, 8, 8, 27, 10, 13, 20, -1, -15, 11, -18, -12, -19, 8, -19, 6, -859, 20, 9, 0, 4, 29, 38, 60, 21, 50, 63, 118, 77, 72, 63, 59, 35, 18, 51, 32, 18, 40, 18, 2, 26, -15, 10, 13, -7, 18, -8, -14, 45, -11, 28, 22, 51, 46, 5, -11, -12, 44, 52, -6, -17, 12, 60, 76, 78, 71, 65, 0, -38, -6, -10, -3, 9, 4, 1, 22, -28, -26, -11, -7, 16, -11, 20, -5, -4, -25, -2, -9, 2, 32, 21, 10, 70, 59, 53, 37, 10, 17, 9, 6, 2, 0, -8, 44, 0, -13, 1, 41, -1, -24, -51, -34, -61, -34, -40, -64, -50, -2, 37, -4, 37, 69, 79, 42, -9, -50, 25, 5, -17, 20, -35, -40, -25, -39, -38, -26, -52, -27, -50, -41, -78, -46, -24, -46, -28, -33, 4, -20, -41, 37, -21, -80, -100, -109, -53, -16, -6, 9, -50, -49, -65, -80, -99, -81, -63, -65, -88, -74, -16, -23, -39, -17, -3, -18, 15, -42, -28, -41, -124, -122, -89, -85, -31, -4, -17, -2, -34, -38, -30, -111, -131, -95, -98, -108, -89, -72, -21, -28, 2, 7, 11, -49, -32, -70, -49, -147, -178, -101, -88, -129, -40, -26, -26, 10, -34, -40, -72, -114, -99, -93, -100, -86, -80, -19, -25, -5, 22, 38, -3, -42, -106, -113, -119, -120, -148, -109, -33, -109, -68, -20, -18, 15, -17, -52, -125, -123, -57, -46, -81, -19, -37, -30, -20, 23, 14, 0, 14, 1, -58, -105, -104, -114, -143, -108, -9, -20, -36, -9, -19, 2, 43, -8, -88, -99, -22, 1, -26, -12, 24, 50, 20, 18, 9, -7, -16, 1, -2, -37, -77, -97, -138, -67, -14, -49, -16, -19, 17, -51, 20, 24, -18, -5, 26, 42, 12, -2, 42, 58, 46, 63, 36, 9, -6, 21, 1, 7, -7, -44, -50, -49, -39, -55, -63, 6, 9, -12, -29, -121, -52, -18, 22, 36, 69, 78, 78, 61, 42, 38, -12, -46, -42, -4, -2, -20, 49, 35, -11, -33, 1, -48, -21, -36, 5, 3, -35, -90, -100, 2, 40, 49, 101, 107, 63, 30, 49, 46, -29, -67, -16, 0, 6, 2, -32, -18, 4, -11, -17, 4, -21, -2, -25, -13, -69, -13, -64, -17, 13, 58, 87, 72, 51, 48, 64, 17, -37, -36, 8, -7, 35, 21, 11, -28, -24, -31, -6, 37, 83, 11, -5, -26, -58, -50, -78, -77, -2, 50, 28, 17, 48, 62, 52, 43, 19, -10, -14, 26, 46, 7, 21, 6, -16, 5, 40, 17, 55, 3, -14, 24, -73, -111, -144, -77, -3, 12, -8, 22, 43, 42, 69, 54, 26, 30, 43, 47, 55, 19, 62, 29, -37, -45, -5, -7, 35, 58, 28, -18, -96, -91, -131, -86, -16, 6, -4, -16, -11, 17, 19, 36, 37, 52, 58, 79, 58, 6, 40, 1, -33, -45, -52, 35, 71, 35, 45, -14, -69, -44, -68, -39, -12, -13, -36, -54, -32, -19, 4, 15, 23, 40, 17, 31, 18, -1, -11, 25, 19, -7, -37, 0, 17, 90, 0, 17, -20, -70, -29, -33, -26, -34, -26, -41, -65, -20, -26, 17, 32, 49, 12, 18, 4, 4, -15, 11, -17, -7, -45, 9, -6, 49, 12, -37, -37, -4, -13, -26, -19, -57, -31, -93, -66, -57, -18, 27, 46, -2, 18, 1, -29, -8, 12, 10, -30, -35, -17, 5, 39, 59, -8, -50, 0, -29, -6, -28, -52, -51, -14, -67, -27, 24, 34, 36, 36, 26, -13, -13, -28, -17, -11, -8, 9, -31, 13, 88, 52, 4, -1, -21, -25, -121, -82, -47, -52, -28, -74, -50, -15, 6, 43, 64, 17, 3, -15, -24, 8, 9, 60, 7, 55, 12, 10, 29, -6, -17, -13, 8, -57, -59, -72, -96, -148, -155, -140, -103, -40, -53, -22, -1, -27, -21, -4, -28, -6, 20, 76, 29, 42, 58, 41, -45, -24, -10, 9, -26, -46, -35, -80, -55, -91, -102, -92, -90, -62, -53, -66, -61, -59, -15, -59, -68, -80, -59, -12, -5, 25, 25, -14, -48, -45, 5, 4, -8, -12, -4, -24, -15, -6, 23, 47, 27, -3, 5, 16, -8, 17, -39, -46, 4, -8, -31, -36, -53, -27, 43, -11, -17, -42, -17, -5, 11, -16, 25, 50, -11, 30, 48, 29, 37, -21, -5, 15, 23, 12, -2, 31, 40, 65, 67, 38, 11, 3, 13, -11, -37, 22, -19, 13, 18, 18, -10, 7, 12, -10, 4, 9, 40, 10, 11, -20, -47, -28, 8, -15, -22, 7, -2, 7, -17, -23, 10, -19, -3, 0, -15, 6, 14, 13, -2, 16, -14, 16, -16, 11, 4, -19, -10, 1, -12, -7, -7, -16, -9, 9, -20, -9, -6, -17, 16, 11, -9, -18, 18, 0, 74, -15, 16, 17, 6, -15, -25, -10, -57, -50, -67, -79, -86, -79, -55, -24, -5, -4, -1, -29, 28, 13, 19, -20, -19, -13, -7, 12, -4, -1, 12, 5, 5, 15, 51, 25, 20, -2, -29, -15, 37, -8, -33, 14, 7, 29, -41, -51, -95, -60, -25, 15, -4, 18, 14, 14, 13, 1, 14, 20, 71, 70, 101, 54, 27, 70, 36, 38, 18, 25, -18, 56, 88, 72, 62, 91, 103, 89, 86, 58, 27, 37, 23, 3, 17, 19, 7, -46, 22, 32, 36, 7, -5, -2, -6, 11, -17, 9, 29, 51, 28, 59, 108, 89, 63, 108, 106, 75, 77, 100, 1, 4, 3, -16, 34, -25, -3, 15, -6, -17, -6, -32, -28, 18, 9, 43, 59, 34, 29, 45, 71, 29, 31, 39, 38, 88, 77, 85, 8, -16, 19, 10, -9, -27, -10, 58, -2, -11, 25, 13, -4, 2, -6, 12, 3, 29, 45, 44, 15, -6, -10, 11, 24, 11, 70, 53, 18, 16, -14, -4, -45, -33, 30, 57, 17, 14, 44, 26, 22, -39, -14, 35, 32, 23, 21, -1, -5, -24, -1, 29, 25, 22, 65, 56, 25, -1, 8, -7, -35, -21, 23, 38, 31, 19, 60, 38, 14, -1, -23, -22, -66, -66, -108, -94, -109, -81, -63, -57, 2, 5, 18, 57, 57, -3, 19, -2, -60, -28, 45, 14, 40, 53, 64, 42, -2, -5, -4, -73, -108, -151, -205, -184, -213, -198, -151, -86, -37, -29, -4, 51, 62, 32, -17, -15, -50, -75, -34, -1, 34, 13, 40, 25, -10, 29, -21, -75, -116, -125, -136, -154, -157, -228, -144, -85, -69, -48, -16, 40, 35, 8, 2, -31, -96, -96, -5, 18, 34, 10, -20, 4, 25, -19, -29, -23, -7, 29, 44, 25, -9, -91, -113, -67, -96, -44, -66, 41, 13, 34, 6, -40, -62, -15, 88, 65, 28, -21, -17, -29, -45, -34, -48, -4, 9, 62, 126, 68, 54, 50, -3, -41, -44, -40, -71, -18, 20, 30, 12, -48, -37, -17, 69, 39, -25, -2, -48, -76, -36, -56, -40, -27, -6, 17, 50, 61, 78, 65, 22, -13, -11, -13, -23, -62, 12, 11, 1, -40, -69, -27, 55, 46, -28, -25, -19, -60, -76, -43, -24, -10, 5, 16, 28, 0, -1, -12, -10, 13, 3, -37, -12, -72, -42, 21, 8, -38, -41, -44, -16, -55, -110, -71, -37, -65, -55, -42, -35, -31, 19, 21, 8, -19, 1, -15, -39, -8, -20, -9, -30, -36, -54, -48, -2, -10, 22, -22, -91, -96, -129, -118, -70, -81, -63, -50, -64, -32, -27, -23, -16, -40, -24, -34, -41, -7, 16, -55, -17, -43, -39, -33, -24, 49, 56, 16, -43, -87, -130, -89, -101, -80, -52, -66, -81, -84, -95, -32, -19, -47, -32, -7, 2, -13, 19, -26, 23, 20, -14, -39, -20, 45, 48, 38, -24, -68, -51, -38, -66, -83, -29, -55, -68, -100, -58, -16, -13, 1, 18, 7, 38, 22, 4, -32, -3, 48, 6, -48, -19, 38, 38, 58, 44, 8, -15, -20, -16, -32, 16, 16, -5, -15, -6, 5, 13, 18, 7, 28, 12, 13, 20, -27, 24, -30, 5, -38, -13, 33, 32, 27, 69, 25, 7, -19, 15, 4, 13, 64, 53, 39, 16, 8, 3, 4, -16, 16, 26, 28, 0, 37, -27, -2, 17, -10, -17, 36, 22, 36, 32, 24, 6, 13, 45, 35, 15, 20, 45, 27, 31, 12, 15, 14, -5, 5, 5, 33, 13, 19, -42, -26, 27, 49, -17, 41, 49, 69, 48, 20, 54, 36, 15, 35, -13, 1, -2, 22, 18, 15, -10, 13, 6, -11, -14, 15, -7, -35, -28, 13, 32, 30, 5, -11, 13, 76, 57, 70, 48, -6, 19, -9, -25, 1, 17, -44, 3, 32, 14, 28, 22, 10, -22, -4, -50, -44, -24, 4, -4, -17, 2, -17, 33, 76, 66, 71, 51, 34, -47, -45, -20, -25, -32, -9, -53, -25, 2, 29, -27, -43, -76, -56, -52, -36, 10, 5, 3, 12, -15, 9, 5, -30, 12, -45, -28, -22, -24, 3, 0, -39, -45, -33, -14, -21, 9, -19, -79, -37, -8, -34, -2, 35, 19, 13, -15, -5, 13, -11, -3, -23, -3, -14, -2, 0, 26, 40, 10, -15, -55, -47, -27, -14, -17, -14, -22, -39, -36, 7, -23, 1, 6, 10, 4, -7, 19, -12, -4, -20, -17, 17, 11, -23, -24, 5, 8, 12, -29, -34, -24, 4, -3, -13, -22, 10, 13, -16, -8, 15, -19, 9, -6, -12, -3, -7, -1, 1, -20, 20, 8, -5, 14, -19, 11, -2, -6, 7, 15, -4, 1, 17, -17, 15, -8, 9, 2, 20, 1, 15, -19, 12, -5, -1237, 2, 17, -6, -14, 31, -8, -17, -10, -12, 13, 33, 33, -32, -3, 62, -22, -41, -11, 11, 2, 3, 17, 25, -4, 3, -20, 7, 5, -11, -19, 6, 22, 15, -49, -70, -41, -50, -72, -87, -135, -154, -161, -113, -123, -88, -105, -78, -6, -44, -18, -50, -60, -8, -5, -16, 16, 6, 25, -31, -40, -24, -15, -2, -12, -15, -2, 1, -40, -47, -22, -43, -68, -63, -99, -102, -81, -69, -57, -73, -46, 33, -25, 12, 18, -10, 25, 18, 22, -29, 23, 4, 35, 103, 38, 11, 10, 22, 40, 29, 27, 5, -63, -50, -120, -115, -86, -101, -116, -47, -5, -10, -18, 17, 48, 22, -2, 16, 9, 11, 39, 80, 58, 54, 44, 30, 27, 50, 57, 12, -37, -14, -36, -74, -48, -71, -61, -62, -38, -7, 3, -19, 34, 21, -12, -28, -11, 13, -7, 50, 72, 43, 35, 45, 47, 45, 12, -2, -16, 2, -46, -35, -7, -31, -51, -60, 7, -21, 12, -8, 16, 6, -48, -24, -41, 17, 21, 27, 32, 46, 27, 29, 42, 48, 43, 61, 20, -6, -56, -52, -52, -100, -105, -72, -20, -8, 23, 10, -4, -58, -67, -60, -85, -42, -18, 10, -1, 45, 32, 30, 32, 56, 99, 85, 74, -1, -39, -92, -122, -181, -132, -87, -18, 0, 14, 45, 18, -58, -61, -61, -99, -64, -24, -26, 19, 6, 18, 10, 63, 73, 57, 70, 97, 15, -97, -173, -232, -183, -79, -37, -23, 31, 20, 50, -45, -67, -9, -61, -109, -100, -53, -51, -2, -39, -21, 15, 40, 69, 100, 86, 39, -65, -200, -240, -234, -197, -94, -14, -42, -16, -30, 5, -39, -88, -29, -17, -63, -80, -42, -37, 14, -24, -2, 8, 41, 50, 50, 51, -52, -186, -269, -249, -173, -133, -49, -38, -17, -31, 7, 16, 26, -37, -32, -22, -74, -90, -80, -69, -46, -16, -7, 22, 53, 44, 18, -22, -163, -196, -231, -160, -114, -79, -16, 37, -4, -24, 23, 24, 49, -15, -13, -52, -57, -113, -85, -64, -36, -39, -14, -12, 71, 58, -19, -111, -202, -157, -101, -70, -19, 16, 9, 53, 73, -24, 19, 28, 75, 10, -6, -43, -72, -55, -46, 9, -23, -34, -31, 18, 30, -10, -116, -118, -138, -65, -25, 19, 49, 93, 10, 53, 88, 20, 1, 35, 48, 28, -51, -58, -2, 7, 39, 32, 6, -14, -16, -18, -18, -88, -116, -103, -62, 46, 51, 52, 80, 61, 11, 28, 76, 23, 8, 33, -41, 3, -9, -30, -26, 25, 34, 38, -6, -61, -31, -27, -34, -47, -34, -50, 21, 76, 76, 84, 53, 85, 52, 50, 64, 41, 6, 35, 15, -69, -56, -51, -9, -14, -4, 11, -17, -65, -49, -18, -45, -34, 21, 39, 65, 91, 46, 81, 34, 70, 38, 64, 113, 46, 2, 44, -8, -76, -53, -16, 17, 13, 6, -4, -25, -6, -25, -10, -15, 36, 20, 39, 78, 30, 12, 17, 24, 54, 63, 17, 14, 28, 41, -29, 10, -59, -51, 9, 18, 14, -12, -25, -9, -15, -29, -29, 14, 39, 9, 25, 1, 25, 32, 51, 59, 85, 46, -5, 35, 38, 38, 17, 24, -35, -18, 24, 14, 20, 33, 12, -3, -8, -46, -57, -47, -6, 11, -34, 4, -14, 28, 73, 51, 61, 74, 25, 30, 53, 12, 20, -44, -65, -11, 65, 42, 22, 26, 32, 28, -18, -39, -38, -34, -23, -40, -47, -24, -6, 40, 32, 14, 51, 67, 17, -5, 0, 15, 23, -24, -33, 21, 61, 32, 21, 21, 25, -27, -34, -74, -37, -51, -36, 3, -20, -19, 4, 8, 10, 39, 31, 33, 11, -28, 0, 7, -33, 5, -1, 33, 67, 44, 75, 24, 34, 8, -11, -35, -25, -26, -29, -18, -34, -32, -23, 4, 27, -25, -22, -33, -32, 29, 5, -21, 3, 16, -29, -24, -31, 30, 50, 41, 32, 36, 33, 10, -23, -59, -50, -59, -51, -1, 3, 13, -42, -45, -26, -55, -9, 17, 10, 9, 12, -35, -24, -9, 1, -4, -57, -76, -31, -51, -37, -44, -66, -88, -79, -100, -151, -135, -84, -96, -97, -61, -71, -22, 23, 24, 14, -16, 15, -2, 14, 14, -21, -6, -24, -73, -79, -43, -94, -39, -17, -1, -29, -51, -114, -101, -38, -10, -37, -12, -20, -18, 3, 11, 10, -5, -18, 9, 6, -7, -32, -42, -30, -35, -26, -34, -36, -30, -23, -16, -74, -78, -67, -72, -39, -2, -30, -1, -4, -5, 0, -17, -17, -3, -18, -21, 2, 12, -20, 7, 13, -10, 20, -6, -11, -19, 0, -5, 5, -11, -2, -14, 19, 7, -16, -9, 15, -9, -6, -7, -11, 0, -874, 9, 15, -16, 17, 40, -26, -49, -31, -44, -57, -27, -19, -102, -77, -51, -31, -32, -32, -34, -4, 4, -15, 12, -15, -7, -5, 10, 19, 5, -12, 5, -25, -51, -67, -97, -40, -13, -10, 19, -18, -52, -105, -34, -52, -18, -47, -99, -73, -51, -94, -85, -84, 4, -9, -14, 12, -19, 27, 10, 18, 17, -33, -34, -27, 19, -20, 13, 21, -28, -14, -13, 11, -15, 18, 13, 58, 29, 41, -19, 10, -13, 11, 7, 10, -16, 12, 35, 1, -22, -22, -26, -7, -48, -59, -22, 24, -4, -2, 2, 31, 20, -5, 34, 61, 57, 44, 22, 52, 30, 38, -16, 7, -16, -7, -51, -44, -7, -10, -30, -18, -34, -25, -48, -26, -9, -23, -9, 4, 13, 38, 30, 60, 45, 30, 21, 26, 32, 55, -6, -13, 7, -22, -53, -3, -11, 30, -45, -16, 8, -56, -35, -34, -25, -19, -15, 0, 21, 20, 53, 25, 61, 17, 21, 2, 37, 43, -6, -20, -24, 28, -8, -31, 52, 2, -16, -3, -16, -27, -22, -1, -27, -14, -14, -31, 17, 21, 37, 47, 58, 12, -44, -4, 31, 64, 17, -11, 14, 4, 1, -13, 43, 36, 42, 29, -14, -23, -21, 2, -39, -73, -60, -2, 73, 99, 67, 64, 69, -1, 4, -17, 8, 9, -15, 7, 35, 20, 37, 25, 63, 34, 28, -20, -15, -17, 9, -32, -51, -88, -1, 57, 88, 78, 56, 52, 24, -18, -13, -24, 17, 3, 36, 8, 41, 50, 60, 69, 64, 35, 8, 9, 0, 30, -7, -45, -84, -98, 48, 124, 116, 69, 56, 18, -3, 17, 19, -13, 51, -18, 11, -8, 68, 50, 8, 33, 49, 0, 5, -11, 39, -10, -35, -64, -90, -41, 123, 156, 103, 56, 21, -14, -3, -21, -23, 21, 61, -5, 34, 19, 25, 56, 64, 91, 22, 8, -8, -4, 42, 33, -22, -54, -30, 50, 182, 149, 91, 52, 33, -42, -49, -36, -41, 1, 18, 12, 59, -5, 10, 39, 39, 33, -22, -9, -17, 17, 38, -13, -55, -39, 0, 112, 155, 108, 57, -6, -28, -52, -65, -35, -23, -28, -40, -17, 37, -3, 28, 67, -5, -15, -34, -33, -19, -26, 2, 2, -29, -41, 45, 119, 113, 72, 21, -34, -49, -58, -71, -48, -85, -77, -3, -11, 5, -7, 49, 77, -14, 0, -33, -45, -25, 11, -21, 0, -39, 6, 50, 115, 131, 64, 1, -66, -52, -80, -102, -89, -63, -86, -1, -12, -23, 14, 11, 33, 29, 13, -37, -46, -17, -19, -41, -17, -27, -43, 35, 114, 125, 54, -84, -54, -61, -97, -83, -74, -23, -41, 15, -43, -13, 11, 13, 28, 62, 28, 18, -20, -16, 3, -15, -39, -43, -47, 25, 118, 118, -8, -90, -60, -23, -31, -6, 0, -24, 28, 10, -53, 16, 6, 43, 84, 1, 17, -12, 25, 10, 2, -12, -39, 2, -15, 4, 81, 51, -69, -61, -66, -24, -44, -15, 7, 2, -6, 21, -18, 1, 22, -1, 53, 44, -10, 8, 39, 2, -5, -11, -36, 1, 15, 16, 33, 4, -43, -74, -44, -18, -43, -14, 0, 0, 41, 17, -6, 8, 29, 51, 35, -19, -30, 15, 33, -8, -7, 7, -41, 15, -3, 20, 2, 39, -10, -59, -15, -42, -45, 0, -28, -22, 47, 36, -44, 34, -1, 14, -23, 4, 24, -8, 2, 6, -11, 15, 0, -3, 7, 16, -13, -11, -40, -11, -23, -22, -20, -34, -14, -14, 63, 47, -31, 73, -3, 48, 46, 14, 55, 44, 39, 40, 41, 23, 38, 46, 39, 42, -17, -30, -41, -34, -39, -20, -7, -5, 17, 10, 39, 66, -21, 29, -12, -4, 73, 73, 32, -5, 19, 18, 32, 25, 39, 21, 31, -3, -14, -43, -34, -45, -41, -7, -33, 0, 5, -3, 21, 35, 0, -19, -19, 7, 75, 36, -5, -79, -50, -47, -55, -15, 11, -25, 17, 2, 25, 3, -8, 8, 35, -3, 7, 2, 35, 17, 8, 52, 30, 9, -12, 7, 32, -18, -20, -3, -20, -22, 25, -1, 44, 40, 28, 22, -27, -34, 45, 27, 43, -5, 45, 10, 40, 23, -19, 39, 0, 6, 11, 0, -17, 39, 18, 25, 49, 43, 51, 33, 87, 21, 30, -6, -54, -72, -1, 15, 39, 8, 11, -6, 19, 9, -26, -11, 21, 14, 9, 6, -5, -1, -19, 4, 52, 25, 21, 12, 9, 21, 25, 2, -5, -22, 20, 11, 11, -5, 27, 29, 32, 25, 15, 5, 9, -4, -7, -3, -7, 3, -14, -5, 9, -5, 20, -17, -19, -13, 17, 3, 6, 12, -5, -6, 18, -20, 18, -16, -2, -6, 16, -15, 9, -15, -13, 1401, 2, -1, 0, 7, -15, -31, -26, -29, -52, -31, -64, -26, -23, -76, -46, -19, -25, -15, -50, -48, -36, -35, -7, -3, 21, -13, -2, 4, 9, -12, 17, -8, -2, -20, -19, -62, -44, -42, -21, -31, -58, -79, -44, -17, -36, -125, -134, -127, -134, -58, -24, -7, 7, -5, 5, -12, -1, 18, 32, 15, 37, 9, -6, -17, -28, -2, -9, -6, 26, -38, -48, -74, -61, -73, -117, -106, -95, -76, -66, -13, 33, -6, -12, -3, 14, 1, 22, 20, -14, 26, 0, -14, 15, 4, -27, -30, -4, -23, -24, -20, -36, -43, -55, -55, -58, -44, -15, 9, 42, -21, -20, -7, 17, 9, 30, -16, 16, 11, 17, 2, -8, -32, -23, -42, -19, 1, -39, -22, -37, -24, -24, -5, -34, -19, 17, 51, 65, 26, 19, -14, 0, 32, 27, 30, 46, 30, 42, -12, 3, 8, -25, 0, -5, -24, -9, 21, 26, 16, 5, -7, -11, -21, 6, 51, 5, 24, -19, -14, -15, 16, 20, 11, 37, 58, 42, 10, -32, -1, -21, -32, -20, -24, -1, 58, 66, 37, 57, 26, 29, 58, 55, 53, -2, 3, -15, -3, 3, -22, -38, -25, 2, 36, 31, -3, -8, 14, -4, -11, 14, 20, 9, 63, 57, 39, 40, 19, 25, 78, 113, 27, 28, 11, -8, -15, -15, -36, -31, 31, 40, 12, 12, 18, -13, -11, -12, -2, 29, 39, 19, 33, 49, 41, 5, 31, 30, 122, 131, 68, 28, -3, -29, -19, 7, -49, -10, 63, 53, 3, 18, 19, 6, 30, 5, 27, 14, 49, 26, 35, 9, -8, 13, 32, 53, 101, 115, 44, 11, -30, -26, -50, -6, -23, -3, 31, 75, 34, 47, 50, 36, 55, 45, 43, 32, -25, -11, -15, 14, 0, 0, 17, 36, 94, 95, 38, 31, -8, -8, -8, -31, -2, 53, 84, 80, 54, 70, 72, 36, 20, 51, 13, 22, -46, -24, 22, 21, 11, 8, 29, 15, 65, 51, -3, 44, -32, -32, -19, -30, 13, 47, 63, 61, 71, 78, 46, 15, 17, 24, -12, -36, -48, -44, 18, 36, 33, 60, 79, 67, 47, 70, 39, -6, 43, 1, 0, -33, -68, -25, 64, 59, 34, 20, 23, 1, -11, -22, -10, -44, -72, -55, 33, 25, 33, 43, 63, 59, 52, 9, -47, 2, -16, 14, 13, -46, -51, -33, 30, 50, -8, -26, -59, -43, -46, -44, -35, -78, -68, -40, 17, 10, 42, 8, 12, 33, -12, -16, -92, -49, -28, 28, -1, -37, -39, -36, 17, -25, -48, -71, -106, -80, -82, -77, -32, -50, -94, -1, 9, 5, 20, -13, -21, -9, -39, -62, -65, -16, -9, 13, 17, -22, -29, 19, 74, 23, -49, -64, -87, -69, -64, -52, -9, -57, -73, -61, 3, -13, 12, -4, -12, -27, -18, -33, -33, -43, -24, -39, -17, -39, 38, 95, 130, 24, -10, -10, -49, -53, -44, 6, -15, -45, -67, -54, 8, 4, -6, 11, -8, -8, -29, -34, -20, -18, -69, -8, -2, -18, 13, 57, 71, 20, 25, -11, -20, -32, -36, -21, -7, -58, -47, -17, -10, -26, -54, -43, -16, -27, -17, -17, -29, -76, -30, -28, 0, -36, -18, 60, 72, 45, 29, -8, -24, -41, -51, -43, -9, -27, -51, -24, -19, -26, -37, -15, 16, -17, 17, 14, -44, -49, 22, -33, 17, 1, 34, 42, 35, 30, 49, 17, -36, -31, -23, -1, -24, -19, 10, 10, -19, -23, -42, -26, 22, 17, 13, 61, -11, -48, 14, -22, -13, -12, 34, 12, 49, 53, 79, 34, 26, 1, -26, -15, -18, 2, -26, -48, -24, -24, -33, 19, 28, 19, 8, 27, -9, -34, 46, -12, -3, 26, 8, -43, 26, 67, 56, 58, 57, 31, 42, 61, 49, 28, 26, -6, -43, 10, 37, 20, -6, -43, -43, -53, -36, -20, -15, -3, -16, 16, -48, 5, 27, 18, 24, 60, 27, 37, 63, 78, 36, -14, -2, -22, -26, -5, 14, -22, -13, -26, -30, -69, -23, -47, -24, -18, -18, -4, 24, 18, 9, -41, 10, 29, 41, 28, 11, 24, 20, 1, 6, -10, 13, 76, 78, 50, 63, -10, -10, -10, 19, -20, -10, -5, -3, -15, -2, -42, -44, 30, 49, 54, 67, 57, 29, 60, -19, -8, -33, 12, 32, 55, 54, 65, 78, 32, 45, 23, 18, 1, -16, 6, -15, -11, -19, 20, 10, 5, 8, 40, 32, -3, 6, -17, -32, -70, -41, -9, 43, 8, 27, 8, 7, 9, 20, 15, -11, 6, -15, 6, 12, 4, -17, -18, 15, 9, 17, 5, -13, -17, 15, 3, 12, -17, 15, 4, -2, 20, 2, 7, -15, -14, 14, -16, 5, -15, 14, -14, -15, -884, 2, -12, 19, -12, 13, -41, -33, -65, -32, -24, -57, -6, -9, -91, -9, -13, -5, -25, -34, -34, -36, -24, -10, -15, -7, -7, 1, 11, -3, -17, 19, -7, -26, -2, 0, -13, -34, -31, -59, -59, -32, -83, -89, -73, -78, -74, -71, -91, -57, -47, -60, 7, 13, 17, -7, -3, -3, 12, 2, 34, 74, 66, 38, -9, -16, -30, -56, -102, -43, -32, -9, -1, -36, -8, 1, -2, -7, -34, -68, -52, 5, 31, 19, 18, 20, 43, 13, -20, -14, -3, -25, 11, -10, 14, -22, -34, 7, 3, -42, -22, -29, -10, 46, 31, 2, -14, -20, -42, 12, 11, -9, 9, -6, 46, -35, -73, -26, 0, -25, 11, -16, 3, 23, 19, 3, 0, -3, 17, 7, 28, 23, -5, 15, -1, 36, 64, 18, -4, 0, -16, 8, 51, -12, -36, 14, -22, 15, 65, 41, 59, 54, 14, 0, 1, -27, -24, -1, 9, 30, -1, 18, 46, 63, 87, 15, -63, 4, -2, 2, -19, -1, 7, -2, 21, 63, 67, 65, 97, 57, 56, 69, 53, 2, -16, -29, 3, 36, 29, 51, 68, 29, 79, 12, -20, -2, 16, -5, -15, -46, 26, 10, 49, 44, 71, 94, 99, 53, 83, 56, 18, -29, -51, -32, -30, 10, 36, 18, 21, -21, -4, 30, 6, -46, -1, 8, -67, -7, 47, -27, 11, 36, 68, 57, 27, 38, 50, 80, 46, -5, -104, -110, -95, -22, 12, -3, 11, -18, 37, 35, 28, -44, 23, -4, -77, -45, -4, -15, -40, 11, 33, 25, 23, 6, 10, 41, 64, -10, -103, -131, -105, -63, -43, -49, -54, -41, 62, 75, -63, -13, -38, -55, -43, -127, -23, -57, -29, -1, 14, -9, -24, -34, -15, 33, 32, -44, -69, -94, -70, -52, -77, -98, -84, -54, -21, 21, -62, -25, 8, -26, -27, -64, -26, -83, -39, -8, -37, -59, -51, -57, -19, 9, 45, -11, -57, -71, -37, -14, -44, -140, -111, -77, -56, -5, -51, 4, -5, -21, -26, -82, -81, -119, -63, -40, -17, -27, -45, -92, -44, -35, -20, -33, -37, -90, -36, 20, 4, -73, -61, -76, -56, -34, 42, -26, 21, -19, -23, -96, -137, -152, -102, -55, 17, -21, -43, -36, -15, -18, -24, -47, -57, -71, -18, -5, 11, -26, -44, -5, -32, -41, -60, -28, 30, 5, -37, -106, -175, -201, -161, -35, 2, 20, -24, -39, -42, -35, -29, -38, -26, -3, -31, 19, 1, -13, -28, -24, -72, 10, -64, -14, -10, 31, 21, -58, -197, -203, -182, -139, -49, -34, -27, -58, -26, -51, -40, -6, 17, 29, 7, -4, 6, 2, -38, -45, -62, -27, -44, -32, -20, 16, 63, 15, -127, -124, -212, -177, -116, -72, -63, -26, -33, -33, 9, 38, 29, 18, 14, 17, 4, -17, -36, -47, -50, -92, -62, -18, -29, 43, 79, 50, -39, -96, -74, -86, -95, -70, -80, -63, -56, 17, 21, 41, 44, 11, 0, 43, 39, -16, -64, -86, -110, -108, -72, -27, -4, 25, 108, 114, 79, -14, 12, 10, -26, -26, -29, -62, -39, 8, 41, 43, 26, 23, 0, 40, 59, 26, -31, -77, -146, -119, -107, -15, -16, 5, 94, 84, 45, 50, 62, 41, 10, 10, -5, 2, -21, 4, 45, 51, 12, -6, -9, 46, 53, 3, -11, -37, -153, -97, -82, -23, -30, 11, 106, 94, 36, 64, 42, 54, 53, 9, 25, -12, 15, 14, 45, -8, -11, -31, -6, 12, 15, 4, -52, -19, -133, -111, -57, -20, -9, 16, 94, 110, 58, 19, 4, -8, 21, 37, 2, -24, -14, -4, 13, -3, -16, -8, 23, -21, -17, -61, -48, -23, -48, -69, -24, 10, 20, -21, -1, 38, 14, 44, 12, -7, -9, -4, -18, -30, -5, 44, 1, -12, 10, 11, 48, 22, -56, -78, -41, 16, -22, -64, 27, 9, 10, -55, 10, 28, 13, 30, 36, 4, -6, 22, -10, -29, 26, 19, 14, -16, -45, -8, -44, -35, -51, -38, -31, -16, -28, -26, 6, 6, 2, 18, 14, 19, -15, -69, -22, 0, -37, -27, -19, -13, 11, 27, -32, -37, -118, -166, -77, -48, -109, -113, -68, -64, 4, 26, 3, -4, -3, 6, -7, 13, -35, -3, -22, -6, -12, 26, 39, 16, 77, 62, 36, 7, -76, -60, -60, -75, -53, -34, -17, 15, -11, -15, 4, 16, -16, 0, 1, -5, 3, 7, -17, -19, 4, 10, -4, -24, 21, 37, 57, -31, -23, 0, -1, 2, 26, 25, -2, 14, 18, -3, -5, 20, -14, 8, 9, 15, 5, 14, -6, -16, 7, 14, 3, 19, -13, 6, -10, -13, -7, -18, -5, 2, -5, 3, 11, -19, -20, 19, 20, -18, -10, 386, 3, -18, -9, -4, 59, -3, -21, -36, -52, -27, -65, -69, -95, -129, -48, -39, -51, -46, -38, -49, -21, -49, 5, 0, 4, -6, 17, 20, 16, 1, -1, -12, -22, -80, -64, -112, -144, -145, -120, -126, -135, -192, -120, -82, -91, -158, -155, -143, -119, -113, -86, -49, 14, 17, 7, -11, -2, -10, -48, 8, -19, -14, -55, -55, -64, -19, -53, -55, -37, -32, -16, 9, -21, -84, -86, -62, -95, -73, -93, -56, 9, 8, -6, 1, -5, 18, -15, -50, -44, -43, -9, 3, -16, 14, 17, 7, -7, 40, 32, -11, -14, -49, 0, -54, -50, -58, -37, -13, 7, 36, -11, -1, 16, 42, -1, -71, -81, -55, 13, 45, 49, 40, 44, 35, 20, 33, 19, -13, -35, -6, 19, -4, 28, 26, 41, 95, 66, 60, -10, 20, 0, 23, -33, -8, -52, -49, 41, 26, 43, 61, 58, 67, 44, -1, 1, -20, -14, -35, -17, 15, 45, 23, 37, 66, 54, 56, 3, 3, 16, -5, -50, -66, -36, -19, 2, 48, 29, 63, 45, 47, 34, 7, -30, -49, -50, -50, -31, -7, -3, -22, -57, 24, 21, 48, 34, 12, 6, -3, -99, -138, -94, -68, 4, 31, 27, 32, 51, 46, 26, 8, -27, -56, -66, -85, -83, -79, -73, -100, -128, -94, 3, 5, 20, 19, 10, -28, -58, -96, -145, -64, -1, 51, -9, -17, -1, 23, 38, 38, 25, -46, -108, -105, -93, -98, -138, -111, -122, -42, 10, -10, -5, 13, 5, -25, -47, -71, -114, -37, 46, -7, -52, -22, 3, 19, 9, 45, 30, -14, -60, -114, -104, -84, -72, -56, -54, 2, 2, 3, 17, -26, -23, -55, -92, -89, -63, -32, 28, 7, -57, -41, -36, 30, 12, 63, 5, -59, -111, -85, -60, -66, -39, -14, -6, 17, 24, 8, 4, 18, -60, -86, -78, -66, -35, -12, 44, 0, -14, -24, -19, -4, 29, 65, 36, -44, -95, -87, -33, 27, 47, 37, 21, -3, 69, 54, 7, -5, -8, -48, -103, -63, -2, 6, -13, -9, -20, -16, -34, 16, 45, 53, 17, -27, -35, -10, 47, 53, 92, 78, 95, 40, 65, 69, 13, 26, -26, -62, -104, -34, -63, 8, -5, 8, 28, 26, 26, 9, 48, -9, -21, -2, -41, -8, 37, 38, 54, 92, 113, 22, 21, 41, 31, -1, -31, -97, -98, -60, -47, -34, 12, -1, -2, 15, 22, -9, -10, -57, -42, -8, 11, 17, 59, 47, 59, 91, 64, -21, -15, 17, -11, 23, -18, -58, -67, -50, -65, -35, -36, -19, 14, -24, -23, -17, 7, -34, 8, 27, 38, 27, 58, 39, 33, 60, 35, -35, 6, 14, 14, -13, -42, 33, 8, -27, -21, -52, -53, -48, -21, -8, -3, -10, -24, -37, -42, -5, -4, 31, 22, -7, -24, -19, 33, 30, 34, -10, -16, 18, -5, 45, 69, 29, -23, -15, 13, 0, 21, 18, 7, -21, -30, -106, -83, -47, -9, 21, -8, 11, -11, -32, -22, 33, 22, -42, 27, -6, 3, 84, 121, 41, -2, 27, 57, 51, 19, 32, 8, 5, -77, -82, -58, -23, -16, -20, 2, 17, 20, -32, -19, 21, -27, -13, -29, -3, -13, 63, 112, 15, 6, -9, 18, 33, 22, 29, -36, -23, -84, -80, -71, -11, -23, -37, -19, -28, 23, 14, 1, 10, -12, -37, -23, -5, 10, 88, 31, 44, -6, 29, 4, 42, 11, -1, -24, -74, -65, -103, -91, -78, -44, -20, -35, -8, 39, -3, 70, 70, 1, -54, 5, 0, 27, 43, 44, 79, 81, 25, 13, 1, 34, -25, -66, -61, -79, -113, -118, -58, -64, -28, -6, 12, 30, 74, 87, 50, -6, -29, -12, -15, -22, -25, 48, 68, 85, 63, 13, 35, 41, -8, -25, -28, -37, -60, -69, -58, -39, 30, 42, 23, 81, 95, 77, 29, 57, 8, -16, -8, -27, -15, -18, 21, 18, 67, 96, 109, 104, -22, -71, -22, -37, -46, 2, 8, 23, -10, 11, 54, 38, 3, 51, 39, 8, -1, -20, 9, -1, -9, -13, -73, -44, 46, 66, 57, 22, -42, -75, -104, -90, -77, -61, -62, -33, -56, -27, -23, -69, -28, 16, 18, 3, 25, -17, 17, 13, -19, -15, -13, -28, -11, -7, -7, -23, -1, -5, -56, -73, -107, -84, -84, -68, -72, -47, -39, -34, -20, 8, -20, -30, 7, 10, -10, 5, -14, -2, -6, -21, -52, -28, -14, -22, -25, -8, -29, 7, 3, -39, -46, -42, -43, -31, -33, -44, -44, 13, 10, 3, 1, -12, 1, -16, -6, 8, 12, 6, -6, -16, -20, 20, -14, -12, 0, -5, 16, -21, 10, 0, -7, -14, 8, 8, -20, 6, -12, -16, -2, -11, 6, -2264, 16, -7, 0, 4, 22, -33, -21, -10, -47, -20, -8, -18, -48, -38, -23, -44, -42, 1, -39, -5, -18, -23, -10, 9, -9, -2, -19, 3, -8, 5, -9, -12, 6, -29, -59, 5, -5, -19, 19, -22, -67, -95, -68, -75, -22, 7, -12, 15, -12, -70, -52, -67, -10, -3, 11, 17, -17, 10, -11, -61, -87, -129, -75, -52, 5, -34, -47, -36, -16, -28, -4, -11, -27, 31, 37, 51, 70, 86, 30, 8, -24, -5, 8, 6, 13, 28, 25, -15, -56, -47, -34, -50, -20, -62, -6, 3, -13, 6, -12, 14, -1, 13, -18, 23, 33, 29, 2, 46, 44, 14, -4, -16, -18, 19, -13, -74, -28, -28, -3, -4, 12, 28, 27, 35, 26, -11, -2, 22, 26, 2, 29, 43, 39, -10, -20, 48, 6, 91, -1, -12, -7, -24, -31, -52, -52, 6, 8, 32, 35, 51, 15, -7, 6, 10, -10, -19, -22, 11, 7, 42, 72, 50, 44, 19, 53, 56, -2, -8, -22, -11, -1, -34, 7, 45, -3, 6, 46, 44, -11, -3, -12, -25, -16, -46, -40, 4, 1, 46, 71, 35, 14, 13, 74, 58, 23, -17, 3, 44, 30, -22, 40, -4, 8, 45, 22, 24, -11, -33, -32, -37, -62, -37, -31, 5, 33, 19, 77, 53, 26, 22, 37, -29, -16, 3, 0, 46, 47, -18, 9, 25, 4, -22, -5, 3, -27, -38, -31, -61, -42, -71, -79, 22, 23, 4, 20, 22, 42, 48, 33, -6, -18, 18, 38, 72, 22, 29, 22, 36, 1, -18, -10, -43, -53, -31, -36, -53, -12, -63, -9, 7, 29, 10, -17, 17, 34, 33, 104, 2, 31, 18, 22, 55, 20, 25, -2, 7, -24, -49, -31, -56, -56, -35, -46, 2, 6, 42, 16, 9, 45, 29, 20, 1, 12, 25, 88, 28, 9, -11, 9, 43, 14, 10, -11, -10, -39, -76, -87, -83, -82, -45, -34, 36, 75, 15, -14, 30, 64, -6, -10, 15, -35, -4, 35, 33, 43, 23, 43, 45, 24, -25, -37, -11, -80, -88, -78, -71, -81, -11, 38, 81, 58, 2, -6, -51, -16, 4, -10, -6, -65, -33, -30, 6, -6, -16, 6, 45, 10, -45, -38, -76, -70, -91, -62, -49, -21, -9, 53, 100, 42, -38, -66, -48, -36, -48, -50, -101, -112, -50, -18, -9, -19, -2, 17, 70, 19, -36, -58, -75, -48, -31, -25, -22, 0, 43, 57, 77, 13, -42, -33, -51, -30, -43, -83, -131, -135, -85, -9, 21, 2, -8, 59, 60, 62, -10, -66, -112, -23, 24, 0, 2, 16, 26, 26, 59, 29, -46, -28, -59, -31, -78, -89, -134, -120, -91, -24, 2, -1, -5, 49, 46, 22, -68, -72, -47, -30, 43, 31, 49, 10, -22, 17, 58, 16, -58, -39, -92, -98, -73, -59, -113, -113, -9, 17, -11, -9, -9, 35, 28, -8, -118, -68, 7, 2, 32, 78, 47, 26, -14, -25, 6, -26, -73, -79, -49, -94, -77, -36, 13, -33, -5, 37, 35, -20, 2, 3, 60, 17, -53, 8, 6, -2, 43, 43, 16, 22, 10, 20, 31, -24, -19, -53, -31, -42, -1, 28, 32, 8, 44, 66, 39, -14, 27, 21, 34, -18, -62, -22, 23, 6, 11, 24, 15, -2, 27, 21, 40, 16, 22, -21, 29, -9, -27, 20, 12, -15, 88, 57, -28, 19, -15, -39, 5, -35, -44, -56, -12, 14, -10, 13, 23, 20, 13, 23, 2, 16, 17, -20, 11, 2, 6, -8, -1, 22, 67, 48, -48, 56, -1, -12, -4, 3, -55, -50, -40, -3, 11, -3, -3, 2, 33, 14, -6, 8, 17, -22, -18, 22, -3, 24, 51, 33, 35, 66, -31, 31, -3, -17, -23, 24, -36, -50, -6, -15, 20, 32, 12, 5, 53, 48, 27, 10, 2, 1, -14, 7, 53, 52, 66, 59, 9, 42, 21, -12, -1, -30, 15, 27, -68, -110, -29, -46, -12, -18, 14, 5, 38, 60, 55, 68, 54, 79, 64, 61, 90, 50, 16, 22, 22, 40, 41, -12, -7, 18, -10, -8, 9, -2, 8, -45, -45, -7, 23, 14, 14, 12, 47, 62, 65, 56, 50, 7, 47, 37, 19, 7, -24, 25, 23, -4, -17, 8, 6, 26, 24, -33, -86, -75, -54, -56, -17, -4, 36, 54, 41, 25, 25, -5, 15, 4, -46, -49, -31, -15, -30, 16, 11, 1, 2, 0, -20, 5, 1, -16, -29, -53, -35, -48, -48, 16, 61, 37, 47, -13, -43, -23, -13, -29, -15, -22, -13, 6, 11, -7, -6, -5, 4, 4, 15, -10, -12, -13, -16, 10, -10, 15, 10, 14, -21, 19, 1, 15, 13, 6, 0, 16, 13, -6, -3, -18, 18, -5, -13, 6, -20, -2378, -12, 1, -11, 16, 25, -8, -14, -4, -27, -18, 27, 46, 15, -32, -10, 14, -37, -37, -15, -9, 1, 3, 19, -3, -4, -18, -10, -19, -6, 12, -9, 15, -29, -40, -54, -52, -72, -90, -6, -11, -21, -48, 7, 3, 12, 26, -2, 26, -17, -47, -46, -51, -25, 0, -6, -10, -17, 20, 7, -19, -41, -89, -108, -67, -57, -56, -36, -6, -52, -23, 35, 15, 27, 58, 62, 54, 32, 27, 39, 49, -11, 25, 0, 1, 12, 7, 17, 23, 2, -42, -45, -33, -60, -23, 8, -50, -31, -17, -16, -6, 5, 13, 26, 50, 61, 9, 20, 71, 76, 41, 7, -4, 18, -2, -40, 22, -9, -15, -17, -49, -13, 12, -22, -8, -6, -18, -10, -23, 4, 10, -2, -2, 40, 6, 20, 38, 55, 52, -1, -2, -16, -4, -34, 42, -7, 7, -17, -27, 16, -14, 3, 7, 11, -12, -13, -48, -14, -26, -26, -30, -19, -36, 30, 32, 70, 102, 8, -9, -23, 11, 15, -8, -7, -27, -13, -12, -5, -11, -10, -13, -44, -24, -29, -7, -20, -1, -33, -11, -29, -15, -23, 6, 66, 70, 31, -25, -16, 63, -3, 6, -41, -16, -15, -14, -32, -28, -34, -21, -24, -5, 12, -1, -31, 0, -7, -40, -54, -34, -24, 17, 64, -4, -12, -16, 37, 32, 47, -7, -19, 6, -2, -36, -55, -10, -13, -9, -4, -5, 10, -50, -48, -36, -14, -40, -27, -29, 6, 0, 41, 18, -25, 14, 28, 50, 45, -23, -5, 2, 6, -23, 12, -24, 3, -15, -33, -9, -16, -27, -2, 1, -22, 8, 8, 8, 6, 29, 91, 20, 13, 20, 12, 58, 22, 4, 5, 11, 3, -50, 16, -15, 5, -8, -21, -1, 7, 15, -6, -44, -23, -5, 7, 12, -4, 46, 63, 41, 40, 20, 37, 75, 54, 27, 52, -1, 46, 19, -5, 19, -8, -9, 12, 19, 13, 17, -20, -14, 45, 30, 48, 30, 16, 85, 53, 17, 38, -14, 48, 79, 60, 57, 54, 16, 44, -5, 9, -27, -33, -12, -13, 2, 36, 31, 26, 45, 35, 47, 37, 65, 54, 32, 5, 9, 22, -13, 21, 86, 124, 40, 33, 20, 38, -1, -4, -5, -20, -4, 12, 31, 53, 69, 67, 68, 69, 67, 44, -11, -65, -15, -15, 13, -2, -2, 52, 91, 98, 94, -11, -17, 29, 11, -13, -13, -27, -28, -37, 28, 52, 77, 85, 63, 2, -60, -118, -164, -201, -178, -72, 13, -21, -17, 17, 26, 127, 63, 2, -22, -18, -17, -15, -14, -34, -17, -22, 6, 24, 54, -19, -68, -154, -214, -311, -290, -201, -136, -25, -11, -11, 11, -27, -8, 22, 7, -52, -53, -50, 10, -5, -7, -6, -24, 2, -27, -70, -108, -149, -258, -339, -277, -258, -186, -141, -92, 24, 9, 19, 21, 32, 17, -46, -116, -87, -65, -45, -24, 0, 11, 11, 21, -41, -147, -210, -213, -243, -226, -216, -136, -114, -69, -38, -30, 17, 36, -3, 29, -27, -41, -101, -187, -97, -31, -24, -10, 18, 46, 27, 0, -57, -103, -165, -124, -95, -59, -16, -25, -31, -27, 5, 32, 55, 36, -10, 9, 0, -62, -118, -192, -104, -15, -9, 16, 7, 41, 2, 0, -6, -26, -11, 20, 39, 37, 26, 16, 47, 22, 8, 61, 36, 6, 35, 6, -10, -33, -91, -116, -85, -51, -25, 9, 23, 11, -7, -2, -7, 45, 50, 40, 76, 57, 31, 6, 33, 57, 21, 62, 90, -5, 53, -10, -46, -34, -107, -116, -92, -64, -35, -12, 9, -12, 5, 13, 18, 29, 51, 32, 35, 29, 40, -25, 32, 55, 40, 27, 48, 23, 46, 16, -34, -42, -58, -105, -83, -63, -64, -29, 1, -25, 3, 26, 27, -4, 26, 40, 35, 14, 7, 30, 30, 29, 18, -9, 6, 44, 18, 19, -39, -49, -57, -80, -117, -76, -52, -12, 10, 21, 16, 37, 33, 16, 22, 33, 73, 78, 35, 81, 32, 42, 39, -4, -2, 47, -1, -10, 7, -36, -5, -32, -96, -86, -66, -46, -26, -36, -8, 42, 19, 57, 53, 62, 65, 73, 97, 63, -1, -7, 4, -34, -6, 12, -3, 14, 6, -4, 20, 10, -32, -98, -77, -61, -45, -21, -23, 21, -6, 2, 16, 15, -39, 3, -3, -6, -82, -65, -40, -20, 4, 9, 1, -9, -13, -12, -9, 3, -30, -76, -60, -85, -64, -76, -8, 40, -10, -17, -54, -61, -64, -20, -23, -23, -19, -36, 8, -15, -12, 9, 10, 17, -12, -8, -12, -21, -10, 18, -13, 20, -10, -5, -7, -12, 18, -5, -35, 4, 5, -13, -7, -18, -8, -13, -9, 10, -10, 5, -17, -19, 880, 6, -14, -7, 18, -13, -3, -8, 20, 5, -31, -30, -39, -45, -39, 3, 4, 2, 16, -10, 28, 0, -12, 23, 0, 6, -14, -8, -10, -10, -5, 8, -2, 40, -7, 13, 30, -14, -12, -15, 16, 59, 102, 42, 7, 83, 78, 49, 79, 86, 95, 51, -10, -15, -1, 1, -19, -19, 15, 26, 6, 10, 43, 69, 81, 45, 15, 24, 108, 96, 65, 53, 75, 113, 97, 58, 88, 121, 123, 132, 81, 8, 10, 18, 8, 15, -29, -14, 63, 55, 68, 76, 83, 37, 38, 27, 106, 37, 52, 58, 20, 46, 40, -18, 19, 96, 109, 96, 117, 32, 1, -14, -9, 0, -25, -5, 26, 82, 114, 94, 42, 72, -7, -29, -21, 23, 43, 33, -7, 9, -5, -34, 18, 48, 60, 16, 31, 40, 59, 4, 10, -2, -25, -4, 5, 13, 48, 25, -7, 0, -1, -35, 5, -19, -3, 1, 1, -6, 14, -60, -50, -35, -8, 25, 66, 69, 36, 8, -27, -7, 13, 1, -9, 55, 90, -12, -26, -18, -50, -27, 3, -15, -47, 10, -15, -15, -39, -29, -31, -17, -16, 51, 95, 80, 59, -8, 3, -32, -30, 5, -6, 47, 43, 31, 9, -44, -47, -68, -20, -11, -29, -17, -2, 0, -16, -9, -45, 0, 8, 56, 119, 164, 21, -37, 3, -8, 1, 3, 7, 0, 26, 28, -3, -17, -1, -4, -15, -33, -32, -40, 23, 40, 20, -27, -24, 22, 65, 108, 97, 137, -18, -3, -22, -11, 15, 21, 22, 50, 53, 47, 7, 13, 54, 44, 13, -47, -69, -18, 29, 4, -2, -53, -6, 1, 54, 76, 12, 69, 56, -18, 3, 78, 36, 34, 24, 37, 53, 96, 75, 101, 112, 62, 33, -37, -39, 30, 60, -10, -25, -33, -4, 1, -6, 1, 18, -16, 33, 1, -6, 41, 29, 18, 21, 73, 124, 112, 99, 179, 95, 82, 15, 3, -11, 4, 50, 27, 15, 20, -1, 38, -31, -40, 10, -4, -6, 1, 21, 25, 67, 18, 106, 144, 127, 125, 160, 145, 74, 70, 8, 16, -14, 12, 9, 51, 40, -10, -20, 14, -42, 14, 51, 27, -34, 11, -12, -2, 13, 35, 61, 141, 109, 105, 106, 140, 94, 51, -14, 8, 0, 6, 47, 49, 22, -16, -51, -6, 23, 8, 26, -3, 7, 13, -8, 1, 12, 39, 68, 104, 114, 95, 138, 152, 116, 20, -3, 8, -5, 14, 20, 49, 78, -14, -45, -17, 23, 57, -44, -32, 46, 12, -13, 7, -54, -28, -11, -16, -4, 13, 49, 104, 55, -14, -11, -45, -43, -3, 21, 58, 65, 46, 39, -22, 6, 8, -41, -2, -22, 5, -5, -42, -93, -106, -80, -95, -42, -52, 0, 1, -8, -9, -39, -64, -53, -39, 4, 48, 109, 53, 53, 61, 68, 28, -15, 29, -24, 4, -14, -16, -39, -106, -81, -47, -43, -14, -12, -27, -35, -49, -77, -99, -77, -78, -53, 55, 79, 97, 65, 88, 96, 37, 15, 62, 29, 28, -1, -3, -12, -52, -29, -2, -1, -23, 8, -15, -64, -65, -56, -78, -70, -79, 9, 68, 63, 63, 66, 43, 33, 28, -8, 40, 25, 32, 1, -13, 15, -29, -21, -18, -25, -18, -11, -38, -15, -40, 24, 8, -25, -68, -43, 52, 79, 63, 102, 65, 47, -2, -43, -5, 32, 47, 1, 16, 18, -9, -10, -45, -16, -14, 11, 20, 16, 16, 22, 20, -33, -15, -60, 18, 40, 83, 91, 86, 120, 27, -45, 13, 54, 67, -9, -5, -21, -48, -11, -14, 23, 27, 9, -18, 27, 68, 38, 31, 15, 9, -6, 27, 68, 131, 140, 107, 65, 31, -48, -32, 54, 4, -5, 31, -20, 17, 19, -19, -17, 26, -15, -10, 34, 38, 31, -9, 12, 48, 69, 109, 140, 187, 173, 124, 18, 19, -27, -41, -51, 2, 14, 37, -42, 14, 28, -25, 27, 77, 77, 11, 26, 41, 33, 29, 17, 22, 62, 89, 95, 104, 145, 93, 12, 29, -53, -18, -9, -15, -9, 9, -12, 26, 77, 68, 51, 100, 73, 63, 33, 23, 54, 55, 51, 22, 34, 115, 125, 112, 95, 71, 42, 36, -31, -42, -40, -16, -3, -10, 1, 28, 58, 57, 50, 91, 29, 1, 45, 66, 0, -18, -13, -9, 85, 80, 80, 56, 36, 39, 10, 3, 20, 14, 11, -15, 3, 3, 18, -15, -5, -2, -26, -14, -29, -1, 31, 84, 60, -38, -46, 47, 24, 47, 14, 40, 38, 24, 9, -13, 11, 19, -15, -4, 17, -11, -4, 10, 1, 15, -16, -2, 2, -2, 2, 0, 13, 20, 3, 5, -6, 13, 19, -1, 19, 18, -20, 9, 11, -13, -2, 7, 3, -592, 5, -18, -21, -18, 38, 8, 31, 5, 28, 10, 25, -14, -25, 19, 57, 23, 1, 68, 17, 29, -9, 12, 13, -13, 1, -2, -19, 18, -3, -5, 16, -20, -19, 17, -6, 23, 72, 16, -3, 18, 4, -11, -1, -27, 13, 20, -10, -26, -70, -43, -42, -87, -20, 16, 11, 6, 15, 25, 8, 16, -29, -45, -17, -13, -1, 27, 22, 15, 17, -9, -27, -13, -34, -28, -83, -76, -59, -39, -29, 23, 15, -19, -15, -4, -11, 9, 24, 72, -64, -65, -42, -51, -15, 8, 27, -33, 25, 23, 12, 13, -21, -55, -66, -31, -43, -50, -31, -64, -78, -16, -1, 0, 18, -25, -33, 7, -54, -11, -2, -42, -20, -49, -29, -18, 28, 54, 56, 39, 25, 28, 23, -29, 25, 41, 1, -39, -101, -64, -11, 10, 11, -35, 14, 22, -8, -10, -18, -36, -52, -36, -34, -10, 13, 54, 61, 78, 41, 55, 67, 39, 49, 52, 50, -5, -72, -27, 5, -11, 4, 45, 28, 55, 73, -11, -25, -18, -21, -23, -59, -13, 6, 55, 38, 66, 48, 63, 72, 47, 44, -8, 27, 8, -87, -39, -18, -1, -18, 43, 12, 37, 48, 9, -16, -37, -25, -47, -37, -47, -8, 38, 73, 79, 49, 76, 43, 68, 41, -1, 19, 3, -37, 11, 23, 8, 8, 46, 28, 35, 9, 3, -21, -19, -70, -33, -42, -18, 5, 44, 61, 89, 58, 55, 36, 36, 54, 11, -42, 22, -68, 7, 41, 0, 25, 43, 38, 42, 20, 1, -57, -52, -25, -23, -17, -25, -4, -3, -21, 29, 12, 39, 14, 17, 11, -2, -16, 21, -64, -1, -20, 15, 40, 90, 123, 45, -18, -33, -32, -37, -44, -13, 16, -29, -15, -20, -54, -39, -16, 1, -3, -2, -3, 6, 16, 2, -61, -28, -25, 12, 76, 82, 75, 12, -2, -35, 10, -40, -19, -32, 11, -18, -28, -29, -72, -35, -1, 9, -10, -51, -42, -26, 6, -24, -82, -16, -35, 28, 51, 40, 45, 39, 7, -35, 2, -14, -16, -10, -43, -52, -35, -58, -42, -45, -16, 30, -13, -54, -67, -55, -24, -42, -51, 19, -19, 1, 27, 89, 37, 28, 21, -8, 23, -3, -10, -24, -55, -84, -53, -60, -73, -41, -5, 18, -45, -86, -47, -77, -28, -100, -65, 57, -29, 20, 33, 14, 77, 80, 21, 20, 25, 7, -28, -41, -45, -67, -86, -96, -128, -110, -62, -46, -64, -76, -75, -61, -81, -105, -84, 83, 22, 6, 43, 9, 94, 82, 46, 58, 44, 5, -27, -46, -43, -39, -38, -71, -96, -99, -56, -50, -56, -55, -36, -12, -70, -95, -45, 33, 51, 19, -14, -83, 9, 36, 79, 70, 60, 14, -25, -14, 12, 34, 49, 49, -10, -33, 15, -3, -10, -14, 27, -23, -56, -62, -42, 33, 70, 2, 2, -11, -41, -1, 40, 27, 42, -3, 12, 18, 43, 122, 138, 137, 134, 48, 47, 34, 39, -4, -2, -1, -11, -7, -7, 88, 25, 21, 36, -21, -70, 8, 42, 25, 32, 13, 31, 46, 44, 82, 75, 94, 41, 37, 45, 46, 24, 17, -13, 0, -7, -15, 20, 20, 47, 8, -32, -124, -138, -43, 48, 30, -6, 22, 23, 12, 10, -9, 9, 34, 21, 44, 33, 68, 20, 10, 17, 4, 5, -12, 0, -3, 48, 34, 20, -103, -73, -35, 24, 32, -2, 20, -8, 24, 12, -18, -11, -16, 31, 29, 41, 52, 10, -12, -12, 23, 18, -21, 3, 16, 6, 10, 7, -44, -96, -59, -15, 14, 15, -46, -40, -26, -17, -14, -11, 15, 5, 32, 28, 47, 27, 16, 25, 45, 26, 12, -13, 2, -29, -4, -23, -17, -76, -37, -46, -50, -25, -46, -33, -16, 4, 6, 19, 20, 32, 25, 12, 56, 41, 71, 6, 6, -14, -15, -19, -29, -15, -3, 32, 6, -45, -100, -60, -51, -43, -62, -24, -52, -25, -3, -4, 27, 41, 54, 15, 27, 31, -17, -16, 25, -28, -43, -32, -7, 15, 4, 0, 4, -13, 28, -32, -82, -89, -93, -54, -54, -51, -24, 8, 3, 49, 20, 3, 0, 39, 21, -30, 0, -9, -42, 15, -33, 9, 17, -3, -8, 41, 43, 77, 24, 11, -4, -46, -29, -68, -31, -36, -11, -16, 9, 8, 38, 30, 42, 15, -8, 21, 19, 16, 17, -11, -8, -18, 17, -19, -13, 27, 28, 21, 24, 17, 21, 59, 47, 9, -39, 25, 21, 36, -10, -22, 20, 28, 14, 11, -15, -18, -12, -5, -3, 0, 14, 6, -16, 14, 12, -5, 19, 18, 8, -16, -12, -14, 22, 26, 7, 7, -13, -13, -17, -13, 8, -12, 7, -8, 20, 2, -16, 810, 3, -9, -3, 20, -8, 13, -3, 13, 3, -17, -60, -47, 9, 3, -1, 35, 44, 5, -2, -10, -5, 19, -12, -10, -11, -1, -21, -11, -6, 8, -16, 35, 32, 0, 41, -20, -20, -20, -7, 16, 19, 70, 51, 63, 27, -1, -26, 0, 24, 71, 41, 88, 4, -16, 0, -6, -2, -9, 11, 31, 55, 26, 66, 2, -38, 20, -18, -32, -47, -45, -1, -44, -44, -31, -55, -73, -67, -40, -72, -61, -7, 21, 13, -20, -19, 25, 50, 99, 119, 98, 89, 88, 26, 57, -29, -46, -60, -63, -46, -35, -17, -13, -3, -17, -49, -70, -61, -69, -72, -48, -5, -15, 0, 3, 63, 88, 129, 133, 86, 71, 20, 16, -13, -28, -68, -36, -16, -33, -51, 16, 15, 19, -21, -4, 0, -17, -10, -36, 20, -5, -17, 10, 124, 152, 158, 83, 88, 74, 10, 1, -17, -18, -29, -15, -31, -29, -33, 2, 28, 22, 39, 68, 39, 21, 2, 15, 1, 14, -13, 75, 119, 164, 108, 78, 60, 68, 38, 16, -9, -11, -15, 3, -20, -49, -30, 18, 25, 33, 54, 37, 74, 48, -14, -4, -8, -13, -17, 31, 126, 97, 68, 42, 66, 52, 62, 35, -33, -31, 10, -10, -6, -40, -16, 13, 11, 36, 34, 37, 47, -6, -38, 23, 20, -11, 29, 30, 75, 71, 74, 55, 35, 52, 56, 14, -22, -11, -17, 22, 1, -23, -15, 35, 31, 77, 62, 39, -9, 6, -2, 5, -14, -14, 28, -55, 66, 60, 20, -17, 16, 19, 21, -22, -58, -34, 1, 37, 3, -5, -1, 48, 70, 60, 65, -5, -21, -14, -30, -51, -2, -9, 53, -66, 46, -30, -56, -23, -1, -3, -12, -32, -36, -37, -3, 1, -30, -16, 32, 75, 72, 87, 46, 35, -19, -37, -23, 14, -14, -14, -1, -6, 95, -59, -48, -15, -51, -28, -41, -31, -27, -6, 23, 15, -7, 6, 53, 69, 55, 85, 21, 9, 9, -49, -22, 0, -19, -14, 1, -44, 63, -33, -71, -32, -31, -27, 0, -37, -31, 0, -11, -10, 17, 32, 84, 94, 109, 113, 51, 25, 21, -14, -21, -32, -7, 9, 8, -9, -8, -17, 2, 39, 35, 6, 21, -14, -4, 7, 7, 11, 46, 8, 68, 106, 87, 105, 107, 65, 42, 9, -37, -50, -29, 4, 25, -3, 6, 64, 129, 85, 52, 2, 3, -17, -28, 0, -1, 2, -19, -11, 31, 36, 59, 99, 104, 52, 68, -5, -50, -69, 10, 16, 1, -51, 25, 183, 146, 64, 40, 5, -21, -45, -65, -19, -13, -52, -51, -46, -37, -26, 36, 31, 88, 95, 52, -14, -39, -47, -36, -15, 4, -26, 2, 97, 72, 13, 29, -12, -18, -37, -87, -59, -60, -31, -35, -65, -34, -23, 21, 50, 70, 99, 40, -15, -30, -67, -10, -3, -53, -84, -35, 60, 3, -36, -15, -32, -5, -28, -32, -26, -4, -17, -30, -5, -1, -3, -14, -15, 9, 24, 6, -23, -47, -53, -43, -2, -27, -51, -19, 62, -36, -43, -10, 13, 13, -3, -26, 8, 9, 1, 25, 6, -19, -27, -31, -45, -18, -10, -85, -74, -13, -15, -60, -8, -35, 13, 34, 57, -10, -63, 2, 20, 11, -19, 26, 5, 33, 50, 21, -9, -48, -39, -73, -46, -23, -43, -76, -56, -29, -10, -36, 11, 17, 36, 58, 67, 6, -1, 29, 11, -3, 5, 30, 5, 27, 6, 21, -18, -58, -64, -67, -22, -53, -63, -98, -64, -84, -14, -82, -21, 7, -7, 75, 6, 30, 10, 2, -8, -2, 23, 26, 12, -28, -33, -30, -50, -35, -62, -33, -53, -68, -95, -144, -8, -53, -20, -8, 18, 24, 21, 23, 7, 9, -2, 31, 19, -4, -14, -18, -55, -15, -36, -10, -13, -28, -63, -51, -40, -71, -91, -77, 2, -13, 33, -20, 2, 33, 42, -45, -34, -4, -71, -61, -51, -59, -36, 2, -34, -59, -23, -6, -27, -32, -26, -30, -5, -7, -48, -65, 0, -52, -25, -21, 8, 8, 1, -12, -23, 15, -11, -33, -67, -52, -68, -33, -13, -43, -6, 47, -31, -36, -9, 31, 10, 15, -2, -6, 3, 23, -28, -15, 1, -1, 8, -23, 35, 21, 33, 30, 4, 21, -4, -5, 16, 69, 124, 105, 87, 74, 64, 56, 101, 86, 80, 47, 24, 2, 5, -7, 14, 9, 13, -12, -17, 41, 49, 50, 50, 40, 54, 55, 31, 82, 64, 68, 83, 64, 83, 33, 45, 67, 67, 1, -12, 10, 18, -14, -5, 10, -20, -16, 18, 7, -2, 9, 13, -12, -10, -3, -9, 5, -22, 28, -2, 19, -17, 12, -15, 14, -9, -7, 20, 8, 8, -16, 15, 1093, -11, -11, 15, 17, 50, 24, 35, 35, 47, 36, 123, 58, 0, 49, 70, 21, 20, 63, 85, 61, 64, 24, 28, 13, -18, 4, 8, -17, 17, 7, -7, -14, 19, 19, 7, 64, 62, 38, 18, 24, 68, 125, 39, -7, 8, 38, 53, 64, 31, 40, 7, -38, 21, -4, -1, -5, 5, 0, 20, 19, 46, 45, 55, -10, -38, -40, -13, -16, -21, -30, -47, -37, 21, -26, -13, -24, -23, -12, 55, 75, 14, -38, 10, 11, -18, -30, -17, -48, 18, 1, 23, 20, -56, -55, -33, -80, -89, -85, -55, -68, -34, -23, -46, -10, 28, 19, 89, 26, -12, -6, 15, -5, -20, -16, -18, 17, -52, -27, -10, -32, -56, -61, -83, -72, -60, -50, -65, -63, -61, -52, -57, -68, 14, 28, 14, 10, -59, -50, -1, 21, 19, -11, 9, 40, -39, -64, -59, -66, -88, -89, -81, -69, -87, -92, -97, -91, -83, -46, -94, -72, -42, -44, -74, -49, -84, -44, -13, 5, 0, -72, -17, 31, -68, -84, -69, -83, -48, -99, -119, -65, -116, -114, -128, -78, -88, -114, -135, -142, -158, -134, -96, -94, -150, -58, -20, 13, -6, -15, -6, -30, -87, -104, -122, -108, -65, -77, -79, -84, -107, -75, -70, -73, -47, -49, -63, -73, -140, -117, -101, -101, -110, -87, -8, -6, -16, -13, -37, -92, -110, -87, -34, -33, -4, -55, -61, -45, -29, 9, -4, 31, 52, 23, 38, 14, -21, -63, -30, 2, -60, 2, 6, -3, -19, 56, -15, -90, -67, -9, 17, 29, 19, -8, 0, 42, 64, 93, 65, 92, 96, 89, 70, 75, 28, 10, 15, -4, -76, -7, -2, 50, -50, 8, -7, -29, -2, 32, 36, 36, 28, 51, 62, 67, 69, 56, 50, 52, 68, 71, 90, 83, 89, 60, 50, 15, -42, -59, -18, 20, 16, -30, -47, -10, -14, 15, 41, 46, 44, 56, 66, 56, 48, 10, -34, 9, -1, 3, 37, 106, 100, 76, 65, 68, -18, -58, -9, 5, 7, 27, 21, -20, 13, 64, 49, 37, 68, 86, 79, 51, 40, -23, -47, -34, 10, 33, 20, 34, 69, 78, 50, 79, 42, 27, -4, -17, -3, -3, 21, 21, 19, 32, 37, 78, 75, 36, 45, 31, 43, -3, -49, -1, 2, 20, 21, 47, 29, 29, 39, 24, 59, 74, 49, 0, -51, 26, 20, 15, -31, -4, 3, -2, 4, 23, 18, 16, 20, -4, -50, -30, 16, 37, 3, 10, 46, 49, -10, 24, -28, 52, 50, -19, 26, 54, 62, -29, -4, 39, -15, 18, 18, 44, 11, 60, 48, -4, -31, 4, 12, 23, 3, 49, 42, 4, -20, -7, -14, 77, 52, 23, 32, -31, -35, -77, 12, 33, 11, 38, 7, -6, 8, 44, 46, 11, 8, 46, 43, 17, 25, 10, 25, 32, -14, -48, 4, 76, 60, 48, 30, -1, -6, -85, -59, 0, 22, 3, 19, 19, -16, 18, 18, 23, 47, 41, 51, 0, 26, 2, 36, 10, -24, -27, 29, 48, 45, 22, 3, -9, -44, -80, -40, 24, 5, -8, 35, 60, 3, -11, 13, 38, 22, 35, 57, 35, 18, -6, -6, -28, -49, -22, 14, 31, 84, 8, -20, -37, -6, 5, -14, 14, -12, 9, 10, 23, 7, 19, 6, 4, 1, -2, 20, 10, 8, 19, 28, -13, -3, -23, 18, 28, 56, -27, -45, 0, -15, 1, 4, -43, -12, -9, 11, -5, 51, 5, 14, 5, 13, -3, 3, 5, 10, 2, 37, 48, -6, 18, 54, 47, -5, 9, -52, -30, -25, -14, -47, -18, 1, -46, 2, -3, -9, 10, 8, 11, -10, 16, 12, 2, 46, 59, 36, 70, 58, 14, 15, 0, -3, 0, -45, -63, -35, 18, 32, -1, -16, -53, -25, -20, -46, -55, -51, -48, -32, -32, -42, -44, 34, 43, 9, -10, 44, -15, -19, -44, 3, 5, -60, -56, -16, 73, 65, 84, 45, 26, -17, -57, -63, -112, -105, -122, -122, -106, -106, -154, -155, -130, -89, -93, -30, -11, 32, -8, -19, -6, 15, -30, -35, -43, -65, -5, 15, -1, -35, -117, -100, -111, -101, -149, -185, -175, -117, -109, -140, -99, -93, -46, -73, -2, -33, 7, -8, -6, 13, 12, -10, -32, -97, -115, -144, -147, -275, -256, -145, -97, -114, -89, -100, -116, -172, -90, -108, -132, -76, -46, -13, -42, -8, 6, -3, -8, 8, -19, 2, 16, -18, -24, -39, -57, -55, -107, -92, -72, -110, -36, -111, -85, -66, -77, -54, -60, -65, -23, -16, -1, -16, 0, 19, -16, -8, -11, -3, -1, 1, 6, 0, 9, 3, 17, 10, 12, 15, -14, -16, -32, -16, 13, 1, 14, -9, -11, 7, -8, 1, -9, 11, -2, -149, 10, -14, 10, -2, -26, -19, -29, -30, -43, -33, -8, 2, -5, -71, -9, -23, -34, -35, 8, -22, -25, -25, -22, -4, 13, -8, 1, 11, 20, -5, 8, -43, -17, -1, -39, -40, -8, -24, -67, -50, -88, -80, -93, -83, -62, -56, -54, -52, -24, -68, -57, -29, -4, 3, 19, 20, 4, 11, 19, 9, -23, -29, -43, -68, -100, -112, -101, -123, -129, -162, -109, -76, -82, -95, -151, -99, -81, -67, -92, -27, 10, 1, 3, 10, -16, 26, 56, 8, -101, -15, -43, -92, -114, -150, -182, -182, -206, -255, -216, -166, -176, -158, -144, -123, -73, -62, -71, -79, -42, -9, 11, 7, -2, 20, -34, -16, -30, -16, 4, -37, -53, -99, -177, -136, -102, -90, -70, -21, -43, -42, -24, -50, -74, -56, 4, -62, -43, 24, 3, 9, -9, 1, -17, 19, 1, -20, -3, 16, 24, -31, -80, -115, -90, -62, -27, -27, -38, 32, 13, 11, 3, -15, 38, 33, 21, 8, -12, 15, 6, 26, 11, 33, 69, 5, 28, 37, 38, -4, -16, -46, -53, -29, -20, -20, 1, 17, 18, 35, 46, -7, 47, 29, 16, 27, 2, 24, -23, 17, 15, 57, 44, 45, 21, 62, 42, 66, 29, 24, -6, -8, -30, 2, 4, 22, 31, 28, 59, 4, 4, 37, 21, 20, -55, 9, 51, 21, 52, 33, 100, 63, 49, 46, 50, 62, 75, 51, 36, -6, -25, -3, 14, 21, 45, 38, 50, -3, 2, 18, -5, 27, -43, -1, 72, -22, 91, 86, 47, 37, 42, 47, 44, 78, 55, 51, 2, 2, 15, 28, -14, 15, 20, 68, 34, 35, 27, 30, 49, -21, -3, 7, 30, 14, 87, 6, 0, 19, 55, 49, 48, 60, 40, 21, 23, 18, 19, 8, 36, 33, 11, 39, 13, 19, 33, 19, 2, 8, -50, 13, 44, 89, 111, 20, -5, 27, 36, 1, 26, 35, 38, 10, 16, 76, 30, 38, 26, 23, 10, -16, 13, 13, 24, 12, 38, -7, -24, 14, 57, 50, 48, -5, -26, -11, 6, 4, 20, 11, 2, 29, 20, 57, 91, 45, 32, 38, 15, 6, -9, -18, -9, -6, 25, -30, -45, 4, 66, 88, 34, -22, 14, 5, -16, -14, -13, -21, -19, 12, 29, 74, 71, 56, 33, 38, -2, -22, -11, -29, -72, -23, 33, -54, -68, 38, 48, 69, 19, 41, 27, 8, 22, -4, -20, -14, -31, 3, 54, 62, 76, 27, 6, 15, -22, -51, -64, -80, -71, -66, -73, -56, -26, 23, 38, -17, 40, 13, 28, 45, 33, 5, -14, -22, -28, 7, -23, 21, -19, -36, -1, -35, -17, -52, -89, -68, -18, -5, -136, -32, -43, -10, -19, -78, -7, -4, 7, 40, 48, 23, 42, -13, -48, -17, -52, -70, -80, -61, -62, -55, -40, -24, -28, -35, 28, -5, -59, -76, -17, -9, -13, -27, -58, -56, -5, -23, -15, -14, -43, -39, -24, -36, -43, -45, -40, -62, -27, -27, -21, -24, -21, -32, 20, 14, -25, -34, 1, -18, 7, -16, -92, -93, -74, -38, -66, -43, -42, -47, -52, -85, -42, -21, -72, -19, -16, 1, -33, -41, -66, -74, -23, -15, -13, -44, -29, 15, -21, -43, -76, -101, -123, -98, -114, -68, -92, -115, -88, -103, -71, -65, -36, -22, 13, 16, -26, -45, -59, -34, -57, -54, -117, -8, 46, 3, 28, 1, -12, -19, -161, -106, -95, -97, -100, -58, -59, -63, -34, -25, -57, -17, 3, 7, -25, -44, -42, -62, -73, -43, -110, 14, -15, 10, 32, -8, 15, -44, -113, -91, -47, -67, -57, -44, -46, -45, -27, -19, -30, -16, 4, 18, 4, -68, -43, -22, -47, -23, -51, -22, -17, 17, 50, 18, 16, 5, -25, -53, -49, -15, -24, -9, -13, -4, 14, 8, 13, 24, 5, 33, 16, 38, -12, -3, -5, 15, -28, 56, -10, 2, 35, 29, -14, -22, 28, -18, -27, -11, 19, -5, -14, 0, -27, 4, 22, 9, 33, 70, 46, 59, 10, 44, -7, -26, -50, -44, 3, -18, 15, 34, 3, 22, 30, 48, 38, -27, 0, -22, -26, -23, -17, -13, 44, 19, 29, 41, 50, -8, 23, 22, -16, -7, 10, -2, -2, 16, -17, -18, 56, 85, 78, 51, 66, 73, 32, 19, 16, 22, 71, 66, 49, 89, 94, 107, 132, 90, 64, 38, 51, 10, -11, 2, -7, 20, 12, -18, 7, 1, 6, 58, 48, 44, 40, 77, 59, 53, 48, 0, 18, 1, 22, 42, 38, 36, 42, 24, 12, 16, -11, -8, -6, -4, 7, 13, -13, 8, 18, 2, 19, -16, -2, -4, 1, 4, 10, 17, 2, -3, 5, 12, -12, 10, 8, 2, -18, 16, 10, 16, 10, 16, -86, -9, -14, -3, -19, 55, 36, 17, -8, -3, 26, 63, -5, -30, -22, 72, 44, 30, 52, 54, 21, 39, 16, 22, -1, 17, 2, 8, 0, 8, -4, -10, -27, -8, 57, 8, 17, 87, 22, -29, 46, 34, 22, 6, 25, 15, 18, 23, 20, -7, -21, -25, -45, -15, 4, 8, 3, 0, 0, 18, 44, 43, 54, 22, 18, 42, 22, 8, 51, -14, -7, 23, 47, 50, 24, 77, 115, 85, 48, 14, 58, 29, -21, 13, 20, 15, 16, 7, 8, -20, -1, 4, -26, 10, -5, 40, 23, 22, 34, 47, 23, 25, 54, 80, 50, 74, 49, 33, 104, 50, 6, 3, 9, 6, 36, -13, 17, -15, 8, 5, 13, -3, -4, 10, 24, 50, 35, 20, 35, 44, 44, 32, 14, -8, 22, 35, 68, 23, 17, -3, 13, -2, 16, 0, 21, 34, 39, 6, -6, 28, 23, 25, 42, 60, 52, 32, 55, 56, 0, -4, -24, -27, -22, -7, 22, 43, 3, 20, -2, -14, -26, 24, 34, 56, 27, 12, 7, 3, 38, 27, 68, 63, 72, 55, 49, -14, -8, -19, -12, -44, -36, -59, 11, 44, -18, 8, 15, -9, 6, 2, 12, 41, 17, -5, 0, 33, 8, 56, 44, 26, -40, -44, -62, -51, -57, -47, -30, -56, -76, -69, -6, 36, 47, 20, 0, -28, -26, -6, 34, 7, -24, 20, 35, 32, 26, 52, 31, -14, -103, -159, -129, -110, -119, -89, -90, -78, -103, -60, -25, 44, 69, 51, -10, -18, -39, -38, -34, -14, 39, 59, 36, 50, 58, 28, -35, -71, -93, -144, -140, -117, -102, -124, -108, -95, -110, -105, -76, 5, -15, 27, 29, -31, 8, -12, 29, 29, 63, 56, 26, 36, 22, -44, -83, -67, -31, -78, -32, -39, -14, -51, -58, -64, -97, -81, -69, 20, -2, 43, 0, 26, 8, -58, 80, 94, 66, 49, 45, -8, -41, -88, -53, -19, -32, -12, -10, 3, 13, 2, -12, -21, -78, -75, -83, -33, 53, 29, 11, -3, 7, -24, 88, 88, 69, 43, 23, -28, -32, -49, -36, 0, -27, -5, -21, -32, -22, 0, 18, 8, -38, -36, -31, -24, 20, 9, 8, -13, 9, 20, 107, 70, -2, -19, -33, -49, -64, -72, -60, -29, -7, -30, -45, -84, -32, -4, 31, 28, -16, -32, -40, -32, 72, 13, 33, -38, 20, 23, 53, 22, -34, -67, -55, -70, -55, -25, -46, -84, -41, -77, -52, -41, -23, 9, -4, 22, 32, -7, -50, -44, 41, 7, -8, -6, 60, 31, 12, 23, -1, -63, -46, -61, 1, -29, -67, -85, -80, -87, -53, -2, 35, 35, 35, 62, 66, -8, -34, -24, 64, 21, 18, -3, 78, 67, 37, -9, -34, -39, -48, -14, 21, -6, -73, -93, -113, -39, 40, 43, 70, 24, 27, 47, 56, 24, 30, 32, 96, 52, 11, 39, 69, 70, 16, -40, 11, 30, -5, -22, -8, -36, -86, -85, -26, 84, 114, 112, 90, 61, 65, 51, 24, 28, 27, 29, 59, 36, 28, 56, 23, 99, 70, -4, 14, 9, 22, 18, 7, -11, -40, -27, 69, 119, 126, 83, 44, 34, 57, 35, 31, 5, 42, -32, 10, 44, 22, -9, -31, 27, 59, 15, 4, -1, 44, 5, 3, 11, 1, 9, 71, 63, 46, 25, 19, 2, 2, 41, 17, 24, -10, -8, -18, 51, 8, 20, 15, 12, 13, 6, -11, 4, 27, 21, 19, 30, 11, 15, 6, 2, 22, 25, 33, 14, 2, 9, 37, -5, -9, 44, 1, 52, 11, 7, 4, 25, 28, -1, -6, 45, 3, 20, 23, 2, 23, -1, 2, -5, -26, -17, 2, -5, -8, -30, 32, 56, 36, 56, 16, 19, 4, 27, 13, 41, -9, 0, 21, -3, 4, 3, -19, -17, 3, -49, -26, -5, -36, -21, 18, 0, -3, -8, 11, 86, 4, 28, 11, 14, -20, -27, 45, 46, 42, 15, 18, 6, -53, -27, 0, -64, -35, -23, -37, -6, -2, 8, 42, -14, -6, -6, -1, -3, 27, 48, -3, -16, 15, -10, 22, -23, -3, -51, -64, -23, -17, -35, -56, -21, 0, -5, -4, 15, 55, 22, -9, 24, 12, 12, 26, -14, -27, -12, -11, -6, 4, 17, 13, -13, -22, 28, 12, 15, 0, 40, 16, 6, -21, -23, -70, -111, -99, -92, -28, -45, -39, -17, -28, 3, 21, 15, -19, -2, 16, -19, 19, -6, -5, 1, 11, -3, -10, -19, -1, -2, -12, -5, -21, -34, 12, 14, -7, -8, -10, 14, 15, 20, 6, 7, 8, -9, -9, -7, 2, -2, 12, -12, -6, 4, 7, 6, 18, 9, 5, 13, 19, 20, 3, -7, -12, 5, 0, -18, 4, 2, -5, 8, 9, 1, -18, -1036, -4, -16, -5, 21, 29, -32, -48, -23, -43, -28, -32, 9, 22, -13, -10, -17, -17, -36, -14, -37, -21, 4, 10, -23, 15, -17, 1, 14, -17, 13, -6, -8, -2, 12, 33, -10, 0, -31, -5, 34, 27, -34, -39, -65, -23, -12, -50, -70, -32, 10, -2, 11, -5, 13, 20, -6, -3, -20, 2, 3, 73, 47, 53, 15, -23, -45, -32, -26, -9, 16, 7, -6, -37, 5, 31, 21, 28, 19, -18, -13, 49, 20, 3, 15, 10, 32, -49, -80, -50, 2, -27, -49, -37, -22, -12, -27, -39, -19, -37, -8, -26, 15, 26, -1, 6, 26, -29, -24, 43, -5, -9, -12, 20, 45, -70, -99, -71, -46, -4, 21, -14, 10, 5, 16, 7, -16, 19, 16, 14, 19, 0, -37, -32, -25, 3, 57, 27, 22, -7, 18, -17, 28, -81, -109, 12, 44, 31, 26, 32, 24, 22, -7, 2, 3, -12, -3, -11, 17, 29, -8, 13, -12, 21, 65, -13, -10, -12, 10, 0, -42, -89, 0, -4, 53, 46, 59, 30, 20, -14, -9, 19, 29, 19, 41, 18, 14, 20, 40, 79, 53, 33, 77, 25, -35, -16, 26, 17, -4, -34, 6, 33, 51, 9, 3, 28, 42, 23, 39, 42, 31, 11, 21, 63, 37, 63, 66, 56, 68, 46, 27, 64, -31, 4, -3, -5, 15, 13, 71, 44, 15, -4, 21, -1, -15, -33, 8, 24, 31, 6, -33, -7, 19, 32, 85, 59, 42, 58, 69, 73, 34, -12, -18, -1, 0, -31, 44, 5, -20, -1, 24, 45, -7, 4, -21, 2, 24, -40, -128, -122, -96, -30, -11, 4, 23, 12, 58, 105, 36, 12, -33, -9, -9, -107, 30, 3, 1, -4, -16, 1, 24, -1, -38, -23, -20, -111, -131, -186, -204, -155, -142, -116, -73, -47, 21, 78, -2, 28, 11, 17, 0, -41, 2, -12, 4, 36, 5, 15, -27, -15, -27, -56, -25, -30, -82, -144, -163, -212, -234, -216, -198, -115, -80, 7, 16, 8, -19, -13, 36, -32, -24, -2, 12, 20, -16, -22, -19, -26, -28, -43, -23, 20, -17, -93, -106, -117, -185, -207, -159, -140, -95, -26, -16, 1, -1, -13, -8, -92, -110, -13, -4, 0, -1, -27, -16, -56, -41, -10, 27, -5, -15, -47, -79, -79, -70, -84, -104, -68, -49, -12, -33, -26, 26, -55, -21, -80, -186, -154, -56, 31, 31, 7, -3, -23, -18, -22, 15, 26, 31, 16, 2, -2, -5, -8, -31, -10, -31, 5, -44, -21, 12, 16, 36, -92, -208, -165, -120, -17, 18, 8, -4, -38, -24, -7, 9, 18, 65, 39, 16, 18, 8, 22, 9, -5, -1, -11, -67, -53, -18, 34, 69, -12, -110, -156, -163, -98, -71, -51, -11, -54, -34, -5, 36, 52, 38, -1, 7, 11, 15, -9, -30, -27, 38, 34, -73, -56, -3, 30, 56, 36, -30, -119, -89, -65, -74, -65, -101, -70, -48, 16, 34, 58, 62, 48, 1, 15, 37, 10, -22, -55, 3, 19, -84, -38, -16, 20, 81, 56, 56, -1, 23, -17, -45, -53, -64, -72, -12, 15, 49, 63, 22, 7, -1, -12, 29, 19, -17, -58, -57, -76, -96, -63, -31, 9, 73, 48, 45, 16, 16, 8, 18, -19, -40, -35, -41, 13, 61, 39, 18, -22, -33, -15, -19, -21, -37, -42, -87, -53, -28, -12, -5, 22, 79, 107, 7, 11, 2, 11, 29, -8, -2, 4, 20, -11, 44, -8, 7, -15, -22, 6, -8, -12, -8, -5, -32, -42, -76, 11, 2, 34, 135, 140, 35, 15, 1, -31, -6, -1, -15, 1, 2, -5, -7, 6, 21, 51, 48, 23, 11, 8, 15, 54, -31, -26, -9, 31, -7, -21, 52, 61, 15, 15, -6, -40, -11, -11, -2, -8, 22, 45, 21, 54, 40, 74, 99, 41, -22, -5, 49, 72, 6, 1, 17, -6, -10, -27, 18, 48, 17, -3, -26, 12, -39, -15, 16, -27, 20, 24, 42, 39, 84, 64, 71, 23, -16, -29, 0, 42, 22, 54, 13, 15, -11, -10, -2, -9, 19, -12, -26, -3, 2, -34, -59, -56, -53, 1, -28, 34, 27, -41, 38, 48, 4, -10, -8, -13, -15, 18, 14, -17, -4, -17, -17, 26, -10, 6, -42, -43, -6, 43, 26, -8, 13, -8, -47, 12, -51, -58, -50, -28, -44, -31, -14, 12, -10, -27, -2, -3, -20, -14, 12, -7, -7, 11, 4, -2, -12, -43, -29, -24, 31, 22, 21, -34, -46, -22, -10, -4, -25, -9, -34, 20, 13, 1, 18, -13, 15, 20, 16, 0, -3, -9, 20, 6, -5, 1, 16, 11, -4, 13, -13, 9, 5, 17, 0, 18, 0, -10, -8, 10, -2, 7, -12, 6, 9, 1336, -1, -9, -5, 18, 51, 21, 12, -23, 18, 12, 56, 58, 67, 62, 29, 41, 39, 63, 23, 32, 19, 14, -1, 19, -2, 20, -5, 9, -10, 14, 1, 11, 4, 7, -5, 12, 78, 77, 130, 56, 94, 97, 130, 56, 77, 109, 92, 55, 10, -45, -61, -44, 16, 19, 21, 15, -17, -9, -18, 80, 74, 38, 18, 55, 86, 64, 121, 77, 67, 117, 131, 161, 148, 171, 117, 85, 53, 47, 22, 37, -24, 1, 2, -15, 11, -8, -53, 4, 16, -25, 3, 41, 45, 17, 50, 51, 58, 64, 58, 34, 13, 4, -38, -25, -20, 5, 29, 87, 62, 31, -3, 14, -7, -30, 9, 1, 6, -45, -70, 10, -43, -24, -1, 12, 35, 31, 22, 3, -26, -32, -44, -90, -50, -26, 7, 68, 72, 26, -14, -17, -17, -39, 30, -35, -27, -33, -27, -12, -7, -27, 0, 19, -4, 39, 20, -16, -20, -20, -66, -43, -23, -12, -32, 5, -18, -25, -10, -19, -19, -75, -12, -46, -60, -57, -20, -21, -37, -48, -54, 5, 9, 26, 31, -26, -42, -26, -29, -38, 9, 1, -44, 12, -12, -22, 19, -1, 21, -15, -28, -33, -4, 9, -22, -46, -19, -67, -23, -13, -4, 20, 37, -21, -51, -63, -58, -44, -25, 20, -22, -25, 4, 26, 34, 9, -11, -52, -40, 37, -18, -34, -14, 4, -30, -65, -22, -1, 29, 31, 25, -60, -77, -82, -58, -38, -44, -10, 24, -29, 19, 48, 27, -9, -64, 0, -110, 7, -30, -14, -14, -25, -49, -68, -32, 6, 38, 28, -12, -57, -48, -77, -55, -79, -52, 6, 13, 0, -6, 33, 21, 31, -37, -44, -127, 3, 19, -35, -12, -39, -75, -67, -14, 51, 33, 17, -37, -51, -51, -80, -109, -75, -77, -6, -25, -12, 8, 4, 44, 13, -40, -74, -79, 34, 41, 1, -49, -80, -66, -31, 3, 6, 32, 27, 1, -46, -63, -28, -69, -112, -105, -95, -44, -31, 19, 5, 23, 3, -35, -91, -75, -16, 4, -5, -33, -73, -35, 4, 13, 62, 79, 64, 36, 8, -15, -7, -54, -77, -127, -79, -86, -54, -7, -3, 27, 21, -7, -58, -89, -14, -29, -22, -22, -33, -3, 14, 41, 92, 96, 66, 62, 37, 31, 33, 34, -49, -96, -79, -64, -64, 9, 80, 29, 4, -15, -41, -61, -68, -71, -44, -42, -4, 19, 18, 65, 115, 85, 53, 57, 47, 48, 91, 87, -1, 5, -73, -26, -6, 5, 47, -15, -1, 23, 37, -31, -104, -50, -32, -19, 6, 9, -4, 53, 125, 115, 68, 10, 27, 58, 80, 64, 32, 20, -25, -2, 20, -25, -4, 33, -3, 43, 112, 67, 41, -19, 14, 15, -6, -29, -18, 41, 85, 102, 83, 37, 28, 55, 38, 32, 41, 17, -19, -43, 11, -6, 11, -30, -10, 9, 69, 95, 20, 5, 6, 1, -23, -65, -56, -20, 55, 67, 27, -15, 30, 47, 79, 32, 30, 53, 29, -17, 24, -49, 0, 7, 22, -6, 94, 114, 18, 37, 53, 6, -19, -34, -39, -21, 7, 26, 28, -20, 35, 71, 36, 24, 49, 57, 45, 0, -6, 5, -10, 65, 16, 53, 40, 90, 64, 40, 25, -37, -11, -26, -3, -21, -7, 6, -11, -26, 34, 25, 31, 42, 48, 90, 24, 52, -15, -12, 10, -29, -42, 3, 31, 74, 11, -10, -42, -35, 15, 29, 21, 32, 4, -9, -12, -23, 18, -14, 32, 54, 59, 38, 7, 29, -71, 21, 3, 70, -8, -2, 36, 63, 51, 11, 13, -35, -1, 24, -16, 15, 16, -6, -8, 6, 29, 28, 52, 54, 81, 27, 44, 64, -47, 29, 4, 18, 18, -7, 27, 47, 2, 2, 19, 2, 1, -28, -44, -30, -22, 7, 0, 22, 25, 52, 47, 27, 7, 37, 39, 58, -53, 51, 20, 21, -21, -23, 32, 67, 40, 5, -21, 20, 21, 14, 10, -27, -7, 29, 10, 23, 30, 33, 21, 1, 7, 12, 14, 24, 16, 40, 35, 3, -16, -6, -5, -1, -27, -2, 33, 35, 39, 14, 22, -13, -30, -25, -16, -18, 0, -27, -25, -31, 10, -10, 26, 9, 41, 23, 35, -11, -8, 9, -7, -9, -18, -3, -29, -21, 11, 37, 33, -18, -27, -16, -96, -69, -142, -153, -95, -97, -61, -73, -43, -20, -10, 2, 15, 5, -13, 0, -4, 1, -2, -35, -19, -40, -32, -59, -53, -59, -32, 14, 19, -80, -66, -23, -26, 1, -42, -16, -37, 0, -11, 10, 20, -11, 14, 15, 19, 9, 17, -5, 12, -10, -5, -6, 0, 6, 17, -10, -2, -10, 11, 0, -20, -6, -4, -20, 11, 0, 11, -6, 0, 0, -10, 2187, -14, -8, 15, 11, 26, 1, -8, 41, 19, 15, 23, -1, 10, 4, 32, 13, -4, -26, -35, -42, -21, -25, 27, -10, 19, 19, -15, 7, 2, 5, 9, -20, 16, -20, 28, 49, 36, 104, 100, 53, 77, 66, 75, 115, 122, 112, 126, 67, 34, 23, 34, 53, 10, 11, 18, -3, -3, 15, -16, -19, 4, -25, 64, 52, 108, 143, 170, 171, 135, 122, 100, 90, 93, 73, 27, -47, 2, -15, -18, 19, 31, -28, 19, -2, 10, -24, 2, 31, 62, 98, 128, 149, 89, 65, 38, 57, 16, 27, 12, 12, 28, -14, 7, -17, -34, -30, -16, -24, -69, -1, -11, 0, 21, -29, 9, 25, 102, 128, 154, 101, 71, 25, -4, 0, -8, -20, -36, -13, -45, -8, 9, 20, -22, 0, 14, 38, -10, -63, -9, -8, 4, -55, 24, 78, 86, 97, 110, 53, 71, 74, 20, 20, -48, -25, -13, -15, 9, -15, 12, -6, 18, -5, 2, 42, 29, -20, 0, 11, -25, -12, 16, 25, 79, 104, 55, 46, 18, 37, 11, 2, -27, -9, -29, 4, -19, -41, -15, -13, -4, -1, 14, 39, -39, -14, 14, 10, 11, -19, 2, 0, 110, 48, 27, -6, 25, -2, -7, -29, -2, -59, -48, -37, -37, -19, -47, -31, -18, 1, 14, 29, -24, 43, -58, -15, -22, 0, 35, 46, 57, 38, -4, -5, 5, 2, -1, 6, -3, -60, -57, -44, -27, -1, -56, -19, -9, 39, 55, 9, 43, -11, -31, 16, -1, -1, 17, 58, 71, -15, 23, 13, 30, 45, 25, 11, 4, -7, -4, 20, -5, -12, -31, -40, 23, 38, 6, 2, 15, -15, -25, -39, -23, 3, 46, 17, 21, 11, 21, 4, 10, 62, 25, 12, 40, 34, 39, 65, 40, 32, 18, 16, -20, 6, -38, -32, 1, 5, -11, -10, -17, 36, 99, -34, -5, -1, -12, 17, 31, 10, 47, 50, 71, 60, 39, 36, 50, 59, 8, -6, -31, -6, -60, -48, -6, -40, -37, 10, 40, 15, 45, -33, -65, -12, -32, -14, 3, 21, 23, 10, 66, 49, 14, 33, 21, 36, -6, -14, -50, -37, -101, -40, 66, 1, -25, 9, 21, 32, 46, -52, -50, -27, -47, -41, 2, 2, 41, 60, 48, 17, -18, 20, 10, -9, -27, -47, -52, -57, -73, -21, -2, 27, 10, 8, 63, 41, 66, 9, 6, -15, -42, -24, 19, 6, 35, 39, 18, 6, -13, 27, 11, -18, -60, -41, -83, -62, -65, -21, 6, 10, 14, -23, -18, -1, 68, 41, -3, -24, -20, -15, -11, 18, 9, -11, -36, -28, -1, -4, 6, -54, -53, -36, -45, -21, -5, 27, 18, 43, 19, -16, -53, 0, 65, 10, -40, -63, -69, -73, -6, -8, -47, -40, -23, -26, 15, 25, 19, -4, 52, 47, 20, 27, 89, 59, -2, 19, -17, 13, -5, 25, 48, -7, -44, -77, -62, -73, -44, -31, -42, -62, -38, -41, 10, 67, 77, 55, 64, 75, 97, 91, 78, 80, 13, 25, 5, -17, 27, 45, 108, 23, -21, -50, -44, -64, -62, -63, -66, -65, -82, -39, 58, 112, 147, 77, 90, 81, 93, 69, 82, 45, 16, 6, 19, -10, 4, 60, 130, 80, 24, -8, -51, -95, -63, -62, -68, -65, -66, -14, 84, 106, 132, 101, 92, 103, 78, 66, 48, 25, 3, 16, -40, -16, 21, 49, 80, 48, -21, 10, -29, -62, -41, -61, -48, -23, -30, -17, 50, 65, 92, 38, 37, 104, 80, 64, 18, -44, -47, 46, -56, -17, 39, 32, 109, 39, 22, -24, -29, -39, -40, -21, 1, 8, 18, 11, 20, 61, 51, 31, 48, 42, 20, 37, -18, -48, -91, 25, -9, -4, 43, 69, 136, 87, 40, 2, 9, -3, -8, -1, 2, -3, -30, 13, 20, 36, 30, -14, 9, 39, 61, -7, -19, -45, -26, 1, -7, 15, 40, 24, 98, 112, 126, 63, 101, 55, -2, -19, 4, -26, -33, -29, -29, -12, -25, 18, 13, 10, 22, 52, 1, -44, -50, -30, -10, -1, -3, 4, 39, 60, 104, 122, 113, -16, -19, -26, -59, -66, -77, -45, -43, -43, -5, 39, 19, 35, 70, 37, 1, 0, -27, -38, 10, 11, 10, 20, -8, 5, 14, 39, 42, -4, -14, -20, 4, -62, -52, 18, -22, 28, 81, 87, 62, 51, 43, 42, 39, -15, -40, -14, -9, 4, 9, -2, -3, 1, 0, 41, 65, 13, 22, 58, -42, -59, -48, -24, -21, -11, -13, 34, 59, 26, 58, 12, 9, 17, -7, -8, -1, 7, -12, -18, 5, -15, -16, 5, 14, -6, 14, -14, 17, -20, 5, -15, 4, 5, 11, 15, -19, 14, -19, 17, 11, -17, 7, -20, 17, 6, 28, -10, 6, 2, -10, 15, 18, 48, 44, 34, 6, 26, 24, 48, 37, 10, -1, 13, 39, 33, 21, 5, 22, 13, -14, 10, -6, -2, 8, -2, 4, 0, -2, 10, 1, 44, 33, 2, 11, 79, 67, 35, 88, 74, 73, 53, 71, 91, 103, 83, 22, -14, -47, -2, -6, -7, -4, 18, -16, -29, -25, 8, -13, 36, 19, -21, 14, 38, 10, 44, 111, 113, 109, 61, 79, 80, 110, 46, 34, 36, 41, -10, -23, 6, 12, 12, -2, -19, -56, 1, 14, 41, 17, 11, -16, -24, -60, -20, -9, 7, 5, 69, 16, -14, -4, -16, -54, -9, -36, -28, -19, 4, -20, 1, 20, -17, -21, 10, 0, -16, 20, 42, 41, 4, 2, -2, 21, 7, 9, 9, -8, -16, -45, 13, -16, -61, -2, -57, -48, -9, 3, 9, -17, 13, 25, -14, 11, -1, 27, -3, 18, -18, -33, -20, -25, -23, -6, -9, -25, -50, -46, -18, 23, 4, -51, -67, -27, -9, -3, -20, -37, 1, 24, -6, -2, 37, -2, -26, -17, -19, -6, -11, -29, -26, -71, -84, -83, -98, -63, -21, -10, -29, -94, -39, -5, 8, -6, 2, -2, 30, 35, 12, -2, -2, -38, -52, -34, 5, 4, -11, -53, -69, -91, -106, -116, -106, -72, -55, -35, -83, -106, -101, -50, -49, -11, 26, 12, 48, 9, -2, -18, -32, -72, -22, -34, -40, -31, -49, -29, -49, -115, -123, -99, -108, -55, -45, -32, -83, -89, -101, -16, -28, -6, 34, 76, -15, 13, -16, -15, -3, -9, -77, -41, -21, -46, -20, 4, 24, -19, -45, -42, -51, -45, -26, -27, -34, -72, -67, 13, -1, 48, -12, 77, -22, 23, -3, -23, -12, -26, -76, -75, -27, 18, 48, 83, 101, 39, 20, -23, -24, -13, -20, -30, -40, -17, -22, -15, 6, 1, 15, 55, -89, -35, -7, -23, -3, -42, -36, -25, 6, 10, 42, 39, 76, 54, 57, 43, 44, 22, 14, -7, -30, -38, 7, -7, 7, -11, 29, 53, -79, -88, -18, -8, -5, -40, -25, -11, 39, 50, -3, 37, 38, 34, 50, 51, 44, 26, -22, 40, 2, -35, 49, -17, -26, -34, 37, 73, -26, -53, -81, -55, -5, 10, -6, -18, 25, 26, 19, 19, 43, 11, 5, 19, 36, 29, 2, 19, -13, 9, 71, 4, -34, -38, 39, 88, 43, -47, -41, -6, 3, 24, -14, -4, -7, -4, 34, 31, -13, -17, -17, 7, 66, 51, 18, 38, 42, 32, 50, 41, -24, 15, 73, 95, 62, -11, 30, 40, 23, 6, 9, -8, -11, -1, 9, 18, 6, -3, -6, 35, 47, 43, 75, 43, 39, 38, 37, 26, -1, 3, 29, 109, 45, 36, 19, 85, 38, 43, -12, 0, -34, -24, 22, 8, 19, 25, 41, 40, 59, 80, 75, 26, 16, 3, 5, 8, -19, 25, 83, 68, -26, -15, 2, 48, 15, 22, 20, -2, -28, 36, 46, 35, 17, 32, 18, 49, 61, 26, 39, 37, -4, -46, -22, -10, 19, 3, 47, 80, -22, -10, 36, 22, 8, -20, -19, 20, 38, 37, 73, 56, 41, 49, 39, 20, 44, 30, 7, 10, -30, -62, -23, -33, -5, 7, 30, 31, 5, 20, 22, 6, -27, -37, -3, 13, 7, 40, 40, 8, 38, 19, -8, 16, 11, 21, 11, -19, -18, -43, 2, -19, 26, -19, -19, 17, -7, -1, 24, -8, -7, 13, -14, -4, -17, 19, -3, 1, -10, 17, -34, -13, -2, -7, -47, -31, -46, -22, 62, -14, 31, -19, 1, 22, 25, 24, 9, 17, -4, 19, 6, -28, 0, -23, -11, -12, -31, -13, -45, -41, -55, -53, -31, -20, -6, -20, 60, -31, 14, 5, -32, -12, 30, 5, 2, 53, -4, -15, -52, -34, -44, -43, -33, -29, -36, -42, -51, -88, -88, -72, 5, -33, -10, -22, 45, 37, -1, 8, -38, 18, 7, -8, -3, 37, 3, -28, 2, -32, -32, -24, -67, -46, -54, -66, -70, -89, -101, -47, -74, -35, -38, -5, 24, 25, 9, -10, 6, -10, -40, -34, -29, -9, -10, -18, -22, -3, -68, -61, -93, -170, -145, -178, -170, -147, -110, -148, -129, -70, -74, -23, -46, 31, -19, 7, -4, -5, -8, -23, -77, -74, -58, -61, -85, -25, -23, -31, -59, -105, -105, -135, -102, -91, -95, -98, -85, -51, -16, -28, -16, 15, 1, -6, -15, -9, -8, -14, -58, -59, -76, -62, -33, -57, -77, -24, 21, 35, -52, -58, -37, -47, -43, -37, -63, -47, 5, -19, -10, -13, -9, -18, -10, 16, -19, -2, -9, -11, 12, -2, 11, 20, -7, 19, 12, 4, 12, 15, 8, -7, -11, -15, -7, -12, -2, -14, 6, -14, 3, 1, -2347, -8, 20, 4, -8, 5, -23, 0, 28, -16, -17, 11, 2, -26, -69, -35, -25, -30, -15, -8, -8, -32, -1, -4, 9, -14, 4, 19, 7, -14, -16, -18, 16, -21, -46, -33, -55, -37, -35, -19, -3, -4, -68, -71, -100, -36, -43, -45, -46, -23, -47, -14, -11, -16, 15, 19, -8, 2, 22, 10, -18, -27, -43, -51, -2, -8, -13, -64, -40, -49, 8, 22, 42, 19, 3, 54, 114, 107, 66, 45, 21, -20, 16, 10, -3, -1, 49, -1, -35, -40, -78, -51, -90, -49, -48, -23, -28, -26, 15, -21, -7, 24, -4, 35, 28, 52, 11, 15, 62, 57, 51, -12, -5, -19, 38, -50, -16, -85, -97, -97, -70, -18, -13, -13, -32, 6, -29, -5, -11, 21, 16, -7, 4, 16, -6, -19, 47, 91, 67, 1, -11, -16, 32, -85, -47, -62, -44, -68, -45, -4, -18, 11, 3, -22, -17, -17, -58, -42, 2, -10, -21, -24, -9, 23, -2, 95, 64, -5, -16, -9, -1, -57, -19, -71, -80, -77, -18, 4, 22, 4, 3, -6, 13, -11, -10, -16, -2, -28, -26, -5, -16, -4, -31, 22, 49, 28, -9, 7, 30, -37, -52, -59, -11, 3, 11, -11, 22, 27, 37, 6, 7, -9, -32, -16, -2, 25, 10, -19, -19, -27, -53, 12, -12, -15, 18, 48, 42, 35, -87, -37, 17, 39, 11, 5, 6, 15, 11, -27, -14, -8, -41, -46, -12, 19, -13, -53, -58, -33, -18, 17, 18, -16, -4, 42, 33, -14, -49, 26, 49, 64, 23, -6, -10, -3, -28, -58, -40, -29, -48, -53, -52, -21, -19, -30, -29, -49, -9, 6, 51, 10, -24, -6, 43, -32, 12, 27, 46, 43, 19, 3, -7, -2, -47, -67, -16, 27, -19, -57, -34, 7, -28, 15, -22, -55, -15, -3, 39, 24, -5, 41, 45, -2, 59, 53, 48, 43, 37, 23, -19, -32, -57, -55, 17, 32, 6, -17, -1, 51, 30, 55, 26, -49, -42, 32, 22, 32, -10, 39, 71, 50, 40, 53, 76, 68, 51, 32, -16, -35, -33, -6, 42, 13, -8, -21, -8, 42, 75, 36, 29, -35, -9, 52, 8, -13, -26, 11, 77, 106, 42, 51, 61, 95, -6, 16, -20, -28, -40, -5, 34, 31, -6, -3, -4, 38, 66, -5, 8, -55, -37, 37, 24, -22, -19, 27, 133, 161, 69, 29, 3, 38, -16, -45, -50, -47, -19, -6, 55, 41, 4, 30, 59, 61, 26, 11, 5, -66, -69, -23, 28, 4, 2, 23, 49, 155, 59, -7, -60, -45, -59, -95, -85, -77, -28, 16, 81, 45, 63, 20, 54, 40, -13, -61, -90, -82, -53, -22, 29, 21, 0, 28, 6, 49, -79, -102, -115, -138, -108, -124, -148, -96, -24, 59, 78, 67, 43, 32, -12, -64, -110, -123, -132, -66, -18, 51, 35, 28, 4, 60, 20, -1, -149, -141, -147, -152, -154, -120, -70, -7, 77, 99, 103, 39, -20, -71, -94, -144, -169, -104, -77, -69, -19, 68, 54, 36, -4, -17, -20, -65, -181, -190, -186, -188, -168, -94, -35, 59, 108, 128, 107, 23, -67, -99, -111, -98, -96, -33, 3, 11, 70, 25, 46, 41, 30, -7, -32, -75, -199, -225, -206, -212, -135, -38, 21, 37, 42, 64, 44, 36, -18, -40, -9, -40, -23, 2, 14, 4, 86, 15, -33, 49, -36, -37, -64, -79, -151, -195, -202, -159, -68, -3, -3, 35, 19, 16, 1, 15, 11, -15, 6, -16, -42, -5, 31, 24, 87, 70, 19, 63, -6, -73, -91, -72, -117, -180, -178, -112, -92, -28, -8, -17, -11, 12, -5, 11, -21, 28, 9, 7, -49, 6, 40, 66, 47, 53, -2, 23, -2, -21, -56, -26, -77, -148, -116, -123, -98, -76, -34, -30, 14, 35, -5, 14, 2, -10, -21, 1, 11, 46, 52, 84, 81, 39, 28, 0, 16, -39, -44, -45, -64, -86, -37, -77, -83, -21, -15, -30, -1, 31, -1, 45, 30, 4, 36, 18, 30, 11, 63, 64, 48, 41, 46, -6, 11, -13, -32, 3, 7, -28, -44, -77, -94, -108, -97, -26, 18, 65, 41, 54, 84, 67, 26, 24, 48, 50, 22, 16, -29, -14, 10, 17, -1, -19, 14, 10, 27, -42, -77, -83, -80, -128, -81, -63, 31, 70, 43, 28, 34, -12, -1, -7, -37, -73, -62, -14, -37, -15, 1, -18, 11, 20, -8, 4, -19, -5, -40, -66, -64, -35, -88, -16, 34, 18, 24, -63, -47, -43, -34, -18, -49, -78, -47, 2, -20, -2, -16, -19, 2, 11, -4, -21, 12, -12, -8, -14, -4, -21, 1, 0, -15, -12, -10, -1, -22, 12, 7, -5, -15, 16, -2, 16, -9, 5, -16, -16, 15, -813, -19, 10, -3, -20, 13, 9, 24, 37, 11, 25, 49, 25, -10, 7, 73, 75, 68, 74, 42, 20, 47, -2, 20, 9, 14, 14, 20, 14, -16, -16, -9, 25, 33, 79, 53, 80, 130, 63, 64, 101, 130, 118, 111, 59, 75, 37, 24, 78, 32, 1, -6, 17, 19, -14, 20, 9, 5, -14, -32, 90, 79, 91, 101, 54, 111, 10, 25, 55, 64, 26, 86, 111, 88, 30, 81, 62, 37, 53, 23, 8, -1, -12, -15, 4, 6, 2, -70, 17, 37, 51, 18, 23, 14, -48, -1, -19, 2, -27, -7, -4, -28, -4, -7, 4, 19, 69, 6, -33, 7, -22, 19, 9, -1, 27, 20, 40, 70, 13, -8, 36, -30, -46, -50, -42, -13, -9, -50, -49, -37, -6, -22, -54, -87, -24, -12, -29, -53, -54, 17, -18, 11, 23, -2, 13, 20, -1, 10, 35, -17, -12, -26, 1, 3, -6, -14, -17, -15, 5, -5, 0, -35, -44, -53, 16, -33, -74, -14, -3, 14, -8, 32, 61, -6, 29, 16, 62, -4, -21, -9, 15, 24, 15, -21, -23, -5, 22, 18, -17, 16, -20, 22, -3, 20, -94, -27, -13, -8, -50, 6, 34, 26, 62, 21, 26, 21, -22, -7, -1, -11, -16, -21, -41, 12, 10, 34, 27, -46, 18, 10, 28, 35, -14, -4, -15, -12, -71, 0, 38, 25, 6, -4, -11, 8, -40, 8, 13, 23, -29, -28, 3, -14, -24, -8, -6, -15, -4, -16, 26, 54, 40, 18, 7, -25, -41, -17, -21, -4, 18, 40, 22, -11, 8, 7, -16, -8, 1, -18, -42, -22, -10, -12, 16, -15, 10, -11, 15, 67, 5, -12, 30, -10, -98, -55, -12, 8, 6, -14, -1, -12, 8, 17, -34, -25, -22, -12, -18, 32, 21, 13, 6, -24, -11, -46, -34, -8, -23, 40, 0, -50, -106, -18, -6, 12, 54, 42, 6, 24, 2, -10, -38, -47, -14, -5, -50, -19, -10, -3, 11, -22, -42, -60, -32, -4, 19, 21, -9, -54, -106, -32, 7, 33, 38, 63, 60, 27, 36, 32, -13, -19, -9, -64, -63, -27, -11, -14, -22, -40, -7, -56, -65, -39, 3, 49, 12, -30, -72, -78, 0, 35, 73, 85, 68, 33, 29, 15, 27, 22, -2, -42, -57, -42, 21, -15, -21, -1, -17, -60, 10, 51, 46, 7, 41, -57, -40, -88, -19, 8, 17, 60, 82, 50, 27, 17, 31, 9, 6, -8, -48, -56, -9, -31, 2, 10, 2, 16, 82, 68, 75, 1, 14, 38, 20, -80, -120, -60, -44, 2, 52, 68, 84, 71, 53, 28, 6, -45, -24, -10, 0, -6, 13, 38, 35, 38, 99, 70, 91, 45, 15, 35, -46, -86, -125, -163, -160, -105, -35, -34, 29, 33, 2, -48, -36, -2, 9, 7, 31, -11, -4, 23, 16, 27, 70, 38, 87, 16, 41, 1, -10, -36, -178, -265, -276, -251, -215, -197, -161, -125, -94, -115, -53, 29, 18, 20, 11, -6, -5, 11, -10, -49, -3, 16, 20, 53, 31, 54, 12, -19, -99, -208, -264, -295, -259, -287, -217, -222, -165, -93, -18, 19, 53, 52, 4, -2, 38, 36, -5, -38, -7, -48, -10, 53, 9, -8, -3, -6, -85, -133, -147, -142, -88, -120, -112, -86, -89, -47, 5, -17, 35, 15, -2, 8, 17, -27, -32, -39, -49, -35, -33, 45, -26, 8, 65, 71, -13, -50, -48, 2, 35, 24, 19, 29, 51, 62, 58, -4, 4, 33, 30, 8, -23, -27, -42, -47, -78, -3, -29, -22, -7, 13, 81, 145, 106, 34, 20, 47, 60, 54, 68, 67, 75, 36, 29, 9, -8, 27, 25, -12, -2, -26, -29, 33, -20, -10, 10, 0, -2, 1, 84, 103, 111, 97, 89, 96, 66, 43, 58, 62, 43, 8, 2, -17, -13, -25, -4, -19, -5, -52, -13, 16, -59, 17, 37, -4, -16, 12, 37, 56, 110, 108, 94, 94, 57, 52, 73, 45, 37, 37, -2, -18, -44, -8, 0, 2, -28, -33, -19, -14, 26, 29, 12, 0, -14, 11, 41, 51, 59, 50, 101, 118, 117, 119, 74, 13, 16, 78, 37, 62, 28, -22, -19, -2, 2, 38, 57, 4, 47, 24, 8, -2, 17, 7, 7, 11, 4, 47, 83, 43, 69, 131, 125, 79, 98, 95, 66, 46, 52, 73, 20, -18, 30, 72, 40, 18, 59, 16, -8, 2, -4, 15, 20, 11, 6, 22, 55, 98, 90, 61, 71, 56, 70, 80, 11, 99, 83, 94, 44, 42, 58, 44, 29, 12, 16, 0, -9, 2, 2, -8, 2, -2, -6, -13, -9, -6, -11, 4, -14, 15, -18, 17, 16, 28, 30, 9, 20, 18, -8, 14, 16, 15, 16, -6, 5, 11, -10, 798, 14, -18, 4, -10, 48, 10, 17, -22, -23, 8, 13, 18, -28, -24, 13, -34, -18, 8, 8, -5, -17, 0, 32, 17, -19, -17, 9, -10, 8, -11, 23, -21, -59, -9, -52, -34, 22, 2, 18, -31, -5, -26, 5, -35, -11, 11, -10, -47, -75, -101, -67, -86, -9, 18, 2, -11, -15, 29, -28, 25, 9, 26, -28, -22, 3, 0, 36, 29, 45, 9, 20, 17, 20, 2, 24, -38, -48, -40, -55, -20, 47, -5, -17, 17, -21, 6, -51, -5, -54, -69, -41, -7, -17, 29, 88, 73, 80, 62, 78, 60, 29, 17, 33, -27, -25, -9, -11, 23, 82, 29, -11, -10, 1, -16, -24, -16, -39, -33, -28, 8, -21, 10, 67, 87, 81, 69, 104, 82, 85, 81, 80, 59, 24, 6, 4, 48, -18, 15, 4, 19, 4, 7, -14, -10, -19, -12, -7, 27, 1, 32, 39, 71, 70, 70, 63, 51, 78, 47, 59, 87, 101, 56, 26, 14, -20, 3, -3, -24, -18, -14, 0, -68, -36, -3, -6, 12, 33, 22, 33, 40, 42, 13, 3, 48, 55, 60, 50, 31, 62, 75, 3, -2, 22, 1, 12, -6, -1, -25, -73, -109, -3, 21, -7, 11, 11, -4, 9, 12, -7, 17, 4, 9, -2, 20, 48, 49, 42, 72, 23, -18, -40, 18, 54, -15, -34, 6, -8, -49, -69, -53, -6, 12, 8, -5, 35, 2, 4, -12, -12, -49, -46, -30, -14, -33, -6, 23, 25, -18, -56, 43, 60, -19, -33, 32, -39, -42, -64, -28, -19, -7, -18, -10, -6, -4, -6, -69, -46, -44, -59, -37, -35, -68, -48, 39, 38, 4, 9, 3, 1, 38, 45, 30, -27, 8, -14, -30, -65, -25, -13, -3, 7, -27, -60, -56, -72, -49, -68, -54, -17, -68, -86, -11, 69, 66, 56, -41, 28, 13, -5, 9, -36, -9, 18, -27, -45, -19, -4, 1, -36, -60, -74, -69, -38, -33, -58, -41, -39, -83, -82, -63, 27, 42, 30, -30, 30, 3, 3, -2, 4, 73, 25, -30, -37, -19, -40, -20, -26, -71, -59, -69, -24, -26, -34, -45, -21, -64, -87, -27, 29, 16, -27, -16, -1, 33, -7, 34, 22, 85, 35, 16, -54, -60, -25, -18, -3, -53, -54, -41, -31, 8, -24, -40, -34, -88, -80, -19, 30, -47, 1, 39, -12, 26, -4, 51, 42, 87, 49, 17, -35, -20, -62, -21, -34, -44, -38, -20, -1, 14, 18, -22, -52, -51, -58, -10, 23, 23, 48, 75, -2, -17, 25, 110, 97, 131, 92, 35, -21, -28, -72, -37, 12, -28, -2, 57, 26, -2, -26, -10, -30, -14, -1, -5, 23, 18, 80, 65, 33, 5, 11, 118, 132, 165, 128, 94, 30, -8, -36, 5, 29, 67, 91, 63, 43, -1, -11, -26, -21, -5, 21, 33, 29, 45, 89, 70, 22, 20, 56, 86, 84, 138, 140, 110, 65, 32, -12, 65, 89, 91, 82, 40, 16, -11, -9, 11, 29, 72, 61, 61, 53, 57, 59, 64, 3, 29, 57, 68, 113, 66, 88, 62, 53, 40, 35, 54, 74, 56, 12, 0, -19, 11, 23, 38, 44, 98, 67, 70, 120, 34, 23, 30, 42, 15, 22, 18, 22, 28, 91, 53, 10, 27, 36, 71, 54, 23, -4, -3, -12, 16, 52, 79, 94, 94, 134, 78, 69, 33, 79, 9, 37, 36, 5, 3, -24, -14, 30, 42, 11, 18, 3, 29, -1, 22, -27, -22, -3, 59, 67, 96, 117, 89, 109, 74, 81, 20, 47, -4, 31, 13, 5, 28, 23, 32, 68, 82, 33, 33, 38, 8, -12, 18, 25, 18, 41, 49, 66, 81, 48, 47, 56, 62, 38, -10, 57, 22, 18, 5, -46, 55, 15, 24, 9, 76, 81, 43, 30, -8, 37, 68, 36, 24, 21, 41, 99, 34, 52, 0, 6, -42, 2, -47, 56, -9, -18, -12, 5, 58, 42, 26, 11, -21, 12, -29, 4, -21, -35, -26, 20, -21, 13, 1, 33, -12, -5, 3, -43, -32, -22, -3, 73, 11, -20, -7, 18, -25, 35, 5, -41, -43, -30, 18, -34, -27, -27, -33, -28, -46, 13, 11, -19, -23, -50, -8, -17, -57, -62, 15, 38, 26, -10, -8, -4, 16, 5, 4, -51, -47, -6, -8, 22, 38, 21, 28, -47, -54, -43, -106, -114, -98, -61, -32, -34, -15, -2, 4, 33, -10, -13, 0, 18, -16, -4, -17, -2, -27, -31, -10, -22, -4, 27, 31, -18, 0, -9, 2, 23, -55, -9, -43, -9, 6, 18, 0, -14, 1, 15, 11, 17, -20, -10, 0, 19, -16, -20, 17, -17, 15, 4, 13, -14, -2, -23, -7, 14, -15, -19, 2, -20, -8, -12, 1, 2, -21, 7, 11, 903, 2, -2, -15, -15, 56, 62, 48, 44, -2, 32, 85, 9, 2, -19, 73, 65, 52, 48, 24, -21, 4, 4, 17, -13, -14, -20, -11, -6, -12, -15, -12, -38, -23, -19, -30, -63, -75, -30, -30, -54, -36, -42, -13, -4, 8, 30, 42, 37, 18, -56, -59, -40, 9, -4, -5, 14, -3, 19, -3, -90, -104, -109, -88, -90, -84, -46, 14, -8, 27, 21, 2, 8, 29, 0, 3, -29, -48, -64, -67, -18, -15, -31, -6, -18, -17, 5, 16, -35, -83, -49, 6, 4, 17, -16, -64, -15, 10, 19, -25, -29, -26, -74, -67, -50, -69, -83, -102, -83, -99, 29, -8, 5, -4, -62, -17, -77, -61, 15, 27, 3, 27, -17, -23, -16, -34, -64, -40, -46, -27, -38, 17, 12, 13, -30, -49, -35, -47, -14, 17, -3, 15, -34, -32, -9, 7, 48, 41, 7, -29, -37, -61, -75, -87, -51, -57, -32, -5, 15, 47, 27, 68, 56, 23, 31, 25, 18, 8, -16, 15, -16, -33, -48, 33, 32, 36, 3, -42, -53, -39, -61, -55, -52, -15, -1, 43, 34, 64, 57, 53, 89, 78, 24, -10, 24, 14, -21, -12, 30, -68, -2, 47, 39, 42, -34, -33, -77, -85, -52, -58, -22, 19, 53, 58, 40, 44, 53, 73, 87, 90, 65, -34, -31, -41, 14, 10, 44, -8, 22, 55, -1, -7, -51, -28, -77, -68, -54, -35, -5, 75, 36, 11, 19, 19, 35, 47, 80, 99, 93, 6, -60, 9, 11, 9, 18, -6, 87, 15, 6, -16, -20, -56, -67, -67, -27, 13, 46, 41, 6, -24, -35, 13, 12, 28, 51, 89, 108, 43, 22, -2, 3, -22, 85, 14, 56, 34, 11, -29, -22, -59, -53, 8, 54, 65, 45, 11, -20, -19, -50, 14, 4, 2, 5, 25, 81, 54, 31, -36, -6, 14, 108, 48, 2, -24, -24, -35, -45, -15, -12, 72, 105, 62, 12, -36, -11, -41, -25, -14, -19, -39, -19, -25, 47, 79, 2, -25, 1, 61, 61, 26, -18, -72, -22, -42, -29, 11, 36, 70, 69, 9, 18, 24, 12, -16, -14, 9, -27, -62, -80, -73, -27, 87, 53, -48, 21, 54, 94, 70, -43, -109, -50, -53, -6, 37, 42, 68, 6, 10, 36, 44, 23, 17, 10, -5, 5, -52, -77, -71, -58, 63, 78, -2, 2, 37, 133, 61, -46, -110, -31, 7, 40, 37, 22, 9, -3, 41, 62, 44, 55, 51, 1, 11, -8, -72, -74, -89, -78, 58, 97, 14, -9, 29, 56, 39, -61, -79, -24, -3, 20, 23, -9, -33, 1, 57, 15, 9, 13, 5, 29, -3, -13, -43, -48, -21, -5, 69, 74, 67, 6, 23, 53, 64, -4, -27, -6, -19, 9, -2, -46, -69, 18, 72, 49, -31, 9, 32, 20, 1, -41, 6, -14, 9, 12, 95, 78, 54, 27, 63, 50, 2, -30, 57, 32, 31, 33, 34, -1, 22, 89, 70, 5, 9, 8, 30, -13, -7, -4, 5, -4, 22, -3, 59, 49, 51, 11, -4, 51, 76, 71, 104, 97, 46, 45, 55, 50, 70, 74, 29, -9, -6, -7, -20, -35, 26, 13, 10, 15, 16, -36, 23, 34, 23, 4, 27, 50, 102, 86, 149, 119, 47, 34, 86, 78, 52, 16, -65, -75, -54, -56, -51, 15, 28, 23, 29, 7, -2, -28, 20, 33, 27, -28, 7, 32, 78, 38, 115, 90, 51, 22, 75, 61, 16, -23, -79, -118, -75, -53, -38, -22, -10, 13, -19, -17, -12, -4, 44, 49, 21, 6, 19, 12, 58, 53, 66, 88, 32, 7, 30, 11, 2, -42, -43, -75, -53, -24, -20, -9, 5, -11, -19, -41, -39, -57, 40, -30, 25, 19, 23, 38, 71, 54, 34, 53, 39, -11, -2, -25, 16, -4, -4, -7, -26, 11, 13, -42, -16, -16, -7, -25, -41, -41, 11, -17, 8, -17, 25, 65, 101, 92, 49, 10, 7, 28, 14, -5, 6, 23, 15, 48, 31, 48, 2, -33, -38, -59, -71, -37, -64, -53, -18, 3, -10, -16, -9, 41, 8, -8, 2, 28, 10, -6, -23, 16, 23, 12, -4, -18, -20, -17, -38, -46, -61, -103, -16, -23, -40, -44, -44, 17, 9, -15, 0, -20, -1, 17, -48, -43, -47, -120, -150, -90, -45, -34, -71, -66, -61, -35, -74, -70, -28, -42, -70, -45, -45, -34, -11, 9, -18, -8, -17, 9, -3, 18, -43, -78, -84, -75, -37, -66, -77, -47, -55, 16, -61, -99, -70, -48, -40, -17, -46, -42, -29, -20, -13, 13, 0, 3, 6, -17, 9, -18, -9, 17, -14, 8, -2, 13, -14, 11, -14, 25, -15, -15, 13, -19, -16, -18, 16, -17, -19, 8, 15, 0, -19, -13, 791, -10, -20, 4, 7, -4, 22, 24, 53, 6, 4, 20, -5, 45, 78, 25, 34, 8, 26, 15, -20, -24, 8, -8, 4, -14, 5, 4, 3, 9, -12, 1, 14, 35, 67, 76, 34, 47, 74, 96, 52, 52, 33, 33, 66, 53, 21, 20, 26, 39, 70, 60, 92, 15, -7, -8, -1, -3, -11, -32, 13, 59, 105, 83, 82, -2, -8, 4, -6, 4, 12, -24, -27, -35, -32, -47, -91, -60, 15, 52, 20, 35, 1, 20, 12, -13, -35, -23, 11, 46, 61, 50, 37, 29, 22, -15, 19, 29, 30, 9, 8, 14, -12, 1, -51, -52, -59, -24, -60, -26, -29, -14, 8, 4, -3, 53, 64, 43, 24, 23, 11, -27, -19, 28, 30, 16, 49, 2, 24, 3, -45, -46, -43, -74, -37, -49, -96, 2, -45, -2, -8, 11, 36, 32, 60, 46, 30, 39, -5, 11, 11, -5, 7, 11, 4, 1, -33, -5, -5, -27, -42, -37, -22, -25, -58, -61, -90, -16, 7, -11, 33, 8, 29, -5, -1, 4, 6, -11, -41, -13, -18, -23, -62, -22, -35, -26, -29, -22, -30, -8, -5, -2, -21, -62, -73, -23, 5, 13, -69, 51, 21, -25, -6, -34, -17, -10, -7, 8, 0, -13, -51, 6, 8, -22, -33, -49, -22, -48, 17, 36, 9, -63, -15, 39, -14, -4, -57, -31, 18, -8, -10, -11, -8, -1, 27, -11, -13, -23, -5, -19, -13, -51, -53, -27, -1, 4, 18, 38, 35, -13, -5, 8, 2, -18, -51, -93, 1, -10, -27, -1, 11, -3, 4, -22, 49, 34, -21, -44, -55, -23, -4, 50, 30, 17, 7, 22, 8, -88, 14, -1, -21, 15, -33, -43, 8, 7, -1, -37, -28, -8, -14, 61, 50, -22, -75, -118, -42, -5, 48, 36, 19, -1, 17, 33, -9, -68, -4, -26, -15, -20, -48, -54, -26, -19, -13, -22, -7, -11, 13, 42, 31, -92, -182, -127, -53, 1, 24, 12, 43, 46, 1, 11, 0, -26, -34, -38, -22, -40, -64, -84, -25, -2, -9, -37, -41, -20, 31, 36, -25, -145, -181, -115, -40, 54, 80, 86, 67, 41, 0, 46, 70, -6, 10, -5, 31, -38, -95, -67, 25, 7, 5, -24, 16, 10, 23, 47, -13, -145, -185, -112, -20, 24, 68, 77, 78, 54, 12, 55, 62, -12, 22, 3, 5, -47, -104, -52, -15, -9, 43, 17, -14, 23, 23, -1, -56, -120, -135, -92, -4, 32, 57, 51, 29, 88, 47, 34, 36, 2, -7, 40, -6, -30, -14, -48, -21, 38, 39, 21, 28, 50, 16, 10, -49, -61, -121, -88, -14, 14, 45, 33, 23, 54, 72, -3, -19, 3, 40, 0, 16, 23, 1, -33, -21, 17, 17, 26, 0, -12, 18, 61, 52, -38, -85, -66, -37, 42, 63, 45, 28, 18, 11, -15, -16, -29, 25, 27, 7, 13, -14, 38, 2, 9, 24, 10, 13, 26, 42, 65, 77, 5, -69, -66, -4, 7, 40, 66, 38, 14, -1, 6, -4, -11, -13, -8, -32, -12, -58, 9, 53, -21, -26, -21, 29, 28, 74, 65, 37, 15, -22, -67, -31, 21, 46, 56, 36, 9, 14, -14, -55, -22, -8, -26, -33, -31, -46, 6, 61, 2, -26, 23, 51, 16, 61, 62, 50, 49, -3, -45, -20, 20, 25, 42, 47, 13, 0, 30, -45, 6, 70, -68, 26, 18, -17, -16, -44, 47, 48, 38, 16, -1, 1, 31, 20, 13, -16, -29, -4, 21, 27, 29, 13, -15, -23, 24, -86, -75, 22, -65, 4, -15, -6, -66, -49, 0, 39, -24, -24, -27, -44, -34, -36, -49, -32, -25, 7, 21, 25, -28, 20, -42, -27, 36, -51, -61, 37, -19, -19, -15, -48, -38, -46, -26, 5, -19, -27, -15, -41, -30, -42, -25, -17, 24, -9, 23, 33, -36, -18, -29, -51, -59, -77, 15, -35, 7, -7, -12, -13, 5, 75, 58, 73, 53, 50, 20, -6, -6, -39, -13, -8, -2, -7, -1, -75, -47, -40, -14, -70, -65, -44, 6, 8, 15, 5, 3, 22, -8, -50, -31, -14, 68, 29, 23, -17, -9, -9, -34, -21, -17, -56, -13, -35, -40, -44, -37, -59, -49, 12, 9, 3, -2, -9, -18, 0, -28, -36, -64, -74, -74, -110, -126, -149, -97, -61, -72, -32, -16, -120, -114, -65, -96, -73, -71, -59, -16, -1, 26, 14, 18, -11, 18, -4, -6, 7, -45, -33, -27, -44, -22, -41, 6, -20, -4, -9, -22, -27, -19, -81, -59, -41, -42, -56, 2, -10, 15, -16, 1, 2, -15, 8, 5, -12, 3, -17, -14, -15, -1, -18, 2, -21, 3, 3, -19, 1, -2, -15, 16, 16, -10, -4, -9, -18, 10, -17, -4, 1, -131, -16, 17, 8, 15, 45, 44, 20, 11, 19, 28, 40, 20, -30, -16, 75, 4, 20, 69, 46, 35, -4, 15, 32, 19, -12, -10, 13, -18, 6, 19, 19, -26, -13, 40, 6, 8, 79, 76, 13, 35, 7, 5, -1, 8, -18, -71, -19, 1, -27, -60, -27, -61, 8, -2, -1, -5, 8, 9, 13, 2, -58, 17, -2, -10, 43, 24, 23, 48, 39, 14, 45, 52, 31, -23, -13, 41, -12, -16, -24, 11, 5, -49, 10, 11, -9, 6, -31, -22, -71, -45, -29, -9, 21, 2, 12, -10, -14, 20, -14, 25, 5, 1, 26, 28, 13, 22, 45, 10, -9, 15, 16, -2, -17, 7, -39, -37, -124, -77, -46, -59, 15, 22, 52, -6, 25, 35, -5, 13, 1, 34, 19, -11, 18, 26, -3, -55, -68, -26, -14, 9, 10, 3, -36, -43, -66, -80, -80, -46, 8, 29, 43, 16, 6, -11, -1, -18, 14, 10, 33, 26, 13, 7, -1, -122, -115, -47, 5, -15, 3, 30, -49, -6, -81, -70, -46, -54, 9, -8, -17, -43, -25, -23, -27, -5, 27, 44, -30, -20, -9, -21, -34, -37, -90, -32, -21, -11, 15, 10, -69, -96, -115, -86, -45, -30, -6, -45, -19, -47, -59, -23, -22, 1, 12, -30, -61, -20, -9, -3, -12, 0, -95, 31, 0, -19, -2, -6, -36, -71, -77, -45, 2, 14, -3, -20, -16, -47, -51, -19, -22, -58, -110, -104, -73, -14, -7, 19, -2, -8, -72, 29, 32, 13, 10, -11, -3, -27, -31, 13, 8, 20, -42, -16, -37, -44, -38, -27, -42, -105, -135, -84, -57, -33, 14, -18, 4, 13, -62, 10, 20, 18, 28, 11, -14, -21, 8, 20, 14, 7, -38, -18, -41, -45, -25, 2, -67, -213, -218, -85, -12, 3, 34, -10, 42, 44, -38, 6, -11, 0, 11, 38, -15, 1, 30, 8, 34, 32, -15, -11, -10, -11, -7, -57, -147, -299, -239, -20, 11, 49, 82, 13, 25, -5, -21, 11, 10, 16, -13, 23, 41, 71, 52, 5, 3, 8, 10, -21, -3, -42, -46, -108, -251, -303, -110, 51, 47, 48, 41, 28, 13, -55, -4, 64, -2, -2, 14, -17, 32, 30, 52, -25, -3, -7, -24, -31, -11, 8, -45, -153, -268, -137, 36, 94, 80, 10, 34, 1, 14, -14, 20, 101, 42, -22, -28, -3, 30, 32, -22, 7, 11, -8, -49, -6, 20, 18, -84, -138, -175, -74, 47, 78, 68, 25, 27, 13, 5, -24, 33, 69, 22, 1, 13, -23, -33, 50, -14, 24, 3, 21, -24, 64, 51, 66, -84, -144, -109, -1, 87, 72, 53, 4, 18, 11, 16, 26, 49, 44, 46, 30, -33, -59, -39, 14, 23, 36, 6, 24, 31, 51, 31, -20, -65, -99, -19, 32, 81, 76, 16, -31, 6, 27, -4, 11, 81, 75, 58, 23, 10, -68, -38, 28, 52, 66, 67, 65, 38, 27, 14, -22, -37, 4, 26, 40, 54, 63, -4, -33, 14, 30, 72, 68, 70, 61, 45, 50, -16, -93, -20, 52, 42, 40, 16, 17, 0, 28, 18, 9, -9, 13, 0, 23, 15, 29, 50, 12, 51, 70, 54, 46, 51, 3, 85, 16, 4, -96, -35, 33, 85, 18, -15, 11, -25, 40, -2, 1, -18, 8, -17, 35, 8, 68, 37, 48, 55, 1, -18, 6, 74, 43, 83, 49, -25, -115, -33, -1, 34, 27, -6, -2, 23, 38, 8, -13, -60, -44, -23, 15, 23, 22, 28, 0, 2, 12, -8, 6, 99, 64, 27, 22, -54, -108, -132, -36, -2, 71, 37, -16, -18, 9, -34, -76, -68, -35, -13, 22, -31, -65, -85, -67, -73, -41, 44, 27, 45, 52, -21, -1, -45, -68, -40, -8, -6, 29, 45, 7, -35, -10, -58, -40, -65, -67, -37, -95, -139, -130, -111, -59, -105, -108, -71, -66, -22, 10, 20, -5, 10, -12, -47, -24, 22, 19, -25, 10, 69, 54, 44, 26, -20, -24, -24, -93, -85, -155, -128, -117, -104, -109, -48, -28, 5, 17, 17, -3, -1, -13, 17, -24, -44, -48, -7, 24, 28, 2, 45, 42, -18, -12, -41, -103, -95, -98, -96, -75, -47, -44, -41, -44, 28, -1, 6, 1, -17, 8, -15, -15, 2, -33, -47, -66, -32, -82, -84, -77, -112, -112, -66, -73, -46, -61, -70, -42, 4, -20, -28, 13, 22, 13, 20, -8, 16, -12, -4, -3, -14, 12, -24, -5, 4, -28, 17, 6, -33, -12, 24, 26, 23, -10, -19, -17, -6, -22, -15, 19, -9, -13, 4, 20, 3, 1, 3, 5, -5, 19, -15, 1, 6, -2, -14, 3, -20, 0, -21, -4, 6, -7, -7, -13, -9, 17, 10, 8, 20, 4, -9, 3, 1232, 5, -9, 18, -17, -22, 7, 49, 16, 14, -34, -44, -32, 25, 17, -54, 4, 15, -41, -16, -7, -1, -6, -44, -2, 7, 9, -2, -14, 9, -14, -10, 1, 40, 42, 48, 28, -2, -24, -2, -18, 7, 41, -27, 32, 12, -39, -4, -13, 16, 51, 39, 79, -1, 0, -8, 9, -1, -14, -1, -8, 1, 24, 87, 59, 25, 56, 76, 47, 2, -10, -33, -93, -68, -52, -66, -74, -52, -16, -27, -22, 8, 30, 14, -10, 16, -9, 21, 32, 33, 73, 81, 109, 98, 152, 70, 63, 6, -29, -24, -7, -33, -9, -25, -22, -58, -60, -51, -53, -75, -43, 14, -13, -8, -69, 15, 36, 61, 84, 114, 98, 71, 65, 54, 40, 9, 8, 7, 1, 0, -26, 14, 10, -15, 2, -30, -70, -27, -61, 13, -19, -8, -2, 31, 18, 45, 67, 89, 62, 50, 69, 28, -7, -20, 7, 33, 9, 10, -3, 35, 7, 7, 44, -13, 0, 38, 8, -2, 2, -14, 39, 10, 26, 48, 35, 58, 51, 44, 10, -18, -1, -34, 11, 6, 8, 36, 3, 30, 0, 7, 20, 10, 5, 2, -36, -9, 8, -17, -44, 6, -3, -2, 19, 13, 9, 25, -35, -22, -37, -31, -18, 8, 27, 6, 30, -9, -10, -29, -8, -2, -33, -48, 8, 19, 5, -15, -55, -37, 9, 47, 0, -15, -46, -51, -71, -51, -50, -43, -51, -18, 8, 23, 5, -13, -18, -18, -10, -43, -51, -79, -34, 3, 7, -16, -84, -15, 2, -15, -27, -53, -68, -69, -70, -57, -50, -34, -21, -24, -2, -2, 27, 17, -4, -9, -30, -51, -8, -51, -57, -8, -14, 34, -81, -39, -11, -43, -14, -73, -72, -70, -82, -50, -25, -53, -44, -70, -1, 13, 40, 28, 21, -3, -24, -24, -14, -20, -16, -16, 14, 4, -43, -12, -69, -10, -27, -84, -67, -53, -33, -18, -20, -32, -45, -83, -27, 31, 42, 33, 48, -8, -5, -26, 9, 0, -39, -9, -12, -24, -66, -13, -26, 9, -23, -19, -36, -22, -24, -16, -30, -25, -53, -8, 8, 46, 54, 32, 54, 37, -1, 5, 27, 10, -51, -35, -4, 6, -21, -15, 1, 26, 66, 29, 65, -2, -35, -18, 3, -10, -18, 4, 12, 37, 45, 44, 77, 69, 93, 59, 36, 16, -46, -4, 11, 9, -76, -41, 55, 113, 143, 77, 40, 41, -27, -39, 9, 23, -1, 5, 23, 24, 29, 60, 105, 143, 104, 94, 72, 11, -43, -20, 20, -4, -53, -15, 170, 134, 155, 104, 54, 24, 15, 28, 4, 10, -4, 22, 5, 20, 65, 102, 91, 129, 121, 75, 51, -5, -12, -20, -10, 18, -22, -20, 114, 71, 99, 70, 50, 5, -1, -8, -1, -10, 19, 15, -7, 53, 66, 90, 69, 31, 60, 1, 30, -27, -31, 19, -28, -23, -82, -84, 21, 50, 9, 30, -3, -3, 4, 3, -30, -36, -13, -31, 29, 13, 17, 29, 29, -5, -19, -14, -4, -14, -48, -13, -39, -43, -47, -33, 80, 62, -47, -48, -27, -12, -1, -2, -37, -47, -23, -24, -33, 1, 6, 34, 3, 12, -42, -14, -49, -28, -52, -55, -29, -11, 4, 7, 56, 21, -39, -16, -63, -10, -9, 24, 5, -35, -16, -9, -35, -19, 2, 27, 25, -16, -20, -31, -61, -23, -54, -27, 49, 39, -9, 53, 29, 7, -3, 16, -21, -15, 12, -4, 50, 43, -14, -26, -28, -17, 19, 17, 6, -3, -21, -52, -66, -107, -16, -60, 18, 30, -37, 9, -43, 4, 37, 26, 11, 8, 1, -8, 9, -2, -27, 9, -8, -3, 10, -35, -3, -30, -20, -117, -102, -85, -6, -16, -4, 12, 48, 15, -8, -8, 22, 48, 5, 26, 2, 2, -22, -4, -1, -2, -18, 8, 3, -18, -25, -65, -50, -111, -37, -69, 12, 6, -12, 58, 33, 1, -1, 43, 28, 10, 6, -21, -20, 22, -17, -1, 4, -18, -22, -45, -21, 1, -24, -40, -61, -55, -7, -66, -12, -20, 19, -19, 39, 39, 50, 43, 22, 9, -60, -49, -11, -24, -24, -33, 28, 21, -52, -23, 4, 12, -4, -23, -15, -3, -26, 10, -38, -2, 11, -10, -17, -23, 22, 39, 58, 87, 46, 10, -4, -24, -16, 23, 34, 29, 28, 35, 46, 50, 90, 118, 83, 36, 37, 15, 21, 11, 20, 13, -3, 11, -11, 27, 38, 59, 88, 80, 89, 45, 50, 63, -2, 54, 101, 82, 84, 57, 46, 57, 44, 29, -5, -5, 6, -3, -9, -10, 18, 17, 6, 9, -13, 10, 17, 3, -9, 12, -13, -17, -22, -3, 18, 13, -4, -18, 0, 8, 16, 6, 21, -11, -9, 9, 1, -1895, 8, 6, -10, -12, 10, -13, 14, -4, 23, 44, 84, 32, 0, 61, 60, 25, 4, 25, 60, 70, 54, 49, 17, 11, 11, 20, -7, 11, -11, 1, 11, 4, 28, 3, -10, 41, 57, 95, 75, 73, 60, 55, 9, 37, 26, 81, 70, 91, 53, -7, -7, -13, 5, -6, 6, 5, -4, 14, 13, -34, -50, -32, -32, -16, 22, 33, -5, 1, -5, 48, 28, 54, 26, 29, 30, 82, 62, 94, 90, 21, -24, 21, -17, 8, 11, 15, -5, -41, -46, -45, -69, -71, -60, -47, -8, -16, -33, 13, 8, -17, -4, -19, -51, -33, 8, 31, 71, 101, 25, 44, 9, -9, -6, 37, -24, -23, -54, -81, -66, -52, -21, 12, 8, -16, -15, 1, -7, -19, 8, -7, -52, -34, -1, -31, -4, 51, 30, 54, 2, -6, -23, -28, -33, -66, -89, -55, -35, -33, -15, -5, -25, -22, -20, 10, 10, -13, -35, -27, -40, -55, -49, -57, -29, 16, 67, 45, 5, -6, -17, -1, -25, -55, -74, -56, -59, -29, -29, -20, -28, -20, 2, 10, 5, -19, -28, -54, -74, -71, -71, -94, -80, -20, 34, 8, 2, -10, 1, 37, 2, -15, -42, -5, 1, 13, 2, -3, 8, 21, -21, 17, 13, -49, -73, -31, -57, -40, -11, -72, -74, -28, 22, -27, -38, -19, 22, 21, -23, -60, -24, -7, 7, 21, 7, 20, 28, 28, 13, 29, -29, -95, -100, -55, -32, -61, -56, -88, -51, -17, -4, 4, 43, 14, 6, 53, 24, -55, -3, 42, 37, 11, 32, 8, 20, 3, -6, 15, -58, -111, -103, -89, -60, -20, -67, -59, -38, -4, 33, 72, 2, 44, 0, 43, 9, -29, 6, 47, 43, 30, 48, 10, 11, 10, -9, 6, -39, -45, -56, -51, -34, -28, -64, -60, -82, -38, 17, 32, 14, 18, 53, 36, -92, 22, 20, 62, 35, 33, 31, 24, 7, -2, -31, 17, -29, -42, -16, 12, 3, -29, -35, -80, -99, -17, 51, 39, 31, -4, 33, 24, -16, 17, 25, 47, 41, 63, 13, 4, 21, -13, 33, -3, -7, -53, -24, -23, -5, -39, -58, -69, -86, -37, 46, 10, 12, -39, 6, 46, 36, 27, 51, 3, 7, 11, 10, -37, -10, -20, 8, 15, -11, -51, -49, -12, 10, -29, -68, -69, -62, 15, 26, 44, -6, -10, 21, 40, 77, 40, -17, 20, -21, -24, -45, 9, 4, -2, -16, 30, -7, -24, -43, 13, -5, -1, -15, -1, -26, 49, 55, 62, 15, 2, 48, 18, 29, -51, -41, 2, -35, -45, -54, -15, 3, -18, 24, 60, 6, -29, -2, 10, -5, 4, -16, -28, 3, 49, 53, 21, 12, 13, 29, 8, -21, -142, -27, -19, -58, -49, -53, -51, -38, -18, 3, 68, 24, 7, 32, 1, 2, -45, -4, -3, 2, 19, 76, 36, 6, 16, 42, -4, -56, -124, -73, -59, -72, -83, -80, -79, -18, 35, 51, 90, 80, 15, -2, -10, -37, -60, 4, 6, 37, 2, 90, 41, 20, 32, 29, -7, -68, -131, -144, -87, -109, -81, -103, -82, 8, 37, 122, 129, 46, 11, -12, -40, -36, -47, -7, -1, 41, 46, 46, 45, 47, 11, 6, -2, -93, -163, -174, -126, -133, -138, -116, -63, 6, 42, 98, 78, 37, 21, -32, -34, -27, -46, -22, -4, -2, 84, 59, 28, 43, -6, -21, -48, -74, -107, -120, -173, -167, -127, -145, -91, -15, -11, 13, 57, 39, 23, -22, -1, -29, -5, 11, 12, 10, 87, 87, 20, 67, 7, -22, -40, -40, -91, -132, -166, -157, -173, -171, -55, -44, -16, -20, 19, 27, 20, 10, -2, 38, -11, 9, 65, 35, 47, 99, 8, 3, 19, 0, -38, -25, -42, -99, -131, -151, -166, -144, -123, -105, -30, -6, 7, 4, 20, 10, 35, 4, 19, 44, 51, 83, 59, 22, 13, 19, -8, 0, 3, -26, -28, -56, -110, -129, -125, -132, -102, -105, -69, -39, 3, 33, 25, 32, 39, 4, 56, 42, 39, 70, 40, 43, 42, 1, 8, -20, -7, 3, 2, -45, -58, -61, -62, -109, -94, -43, -22, -33, 2, 34, 77, 79, 45, 3, 29, 46, 7, 30, -23, 22, 42, -6, -1, 1, 6, -4, -4, -6, -41, -9, -44, -73, -77, -104, -26, -16, -7, -20, -4, -9, 9, -23, -18, -98, -64, -38, -2, -23, 17, -4, 9, 0, 5, 17, -16, 11, -1, -3, -28, -18, -35, -22, -38, 1, 6, -65, -57, -43, -48, -42, -70, -57, -33, 8, 19, 18, 10, 1, 17, -8, -11, -6, 3, -14, -1, -17, 13, -15, -5, -17, 0, -15, 16, -5, -23, 1, 15, 11, 1, -15, -7, 18, 8, 17, -7, 7, -6, 613, -16, 21, -4, 1, 5, -16, -16, -30, 25, -11, -35, -26, -3, -6, -91, -35, -12, -36, -19, -8, 23, 7, -37, -1, 15, -5, 10, 17, 1, -20, 9, -6, 15, 31, 24, 64, 21, 54, 59, 27, 18, 48, 18, -5, 31, 9, 9, -18, -6, 53, 42, 70, -3, 0, -14, 8, 15, -7, -18, 14, 21, 50, 40, 91, 85, 65, 45, 11, 26, 59, 34, 8, -6, 18, 24, -15, -1, 31, -26, -66, -17, 12, -18, -8, -16, -34, -50, -40, 17, -9, -47, 21, 19, -33, -81, -2, 10, 2, 8, -2, 11, -7, -6, -6, 10, -6, -51, -24, 8, 26, 8, 2, 3, -47, -36, -31, -7, -80, -93, -34, -89, -70, -52, -21, -2, 27, 25, 18, -7, -6, -20, 37, 2, 6, 1, 22, 23, -15, -15, 4, 17, -67, 12, -24, -55, -117, -103, -54, -69, -90, -57, -52, -6, 22, -13, 3, 29, -12, 11, 51, 70, 65, 63, 76, -7, -21, 2, 13, -4, -39, -35, -45, -65, -65, -64, -43, -61, -61, -42, -59, -24, 10, 12, -19, -1, -9, 24, 32, 67, 56, 74, 37, 6, 6, 27, 16, -6, 14, -25, -49, -48, -62, -68, -54, -9, -37, -25, -36, 9, -21, -5, -41, -35, -47, -52, -46, -1, 24, 28, -9, -31, -8, 16, -8, -11, -9, -36, -89, -107, -84, -82, -46, -18, 4, -30, -14, -6, -14, -23, -77, -105, -76, -131, -90, -85, -7, -7, -43, -62, -15, -23, 12, -56, 21, -71, -117, -133, -133, -101, -38, -69, -42, -36, -25, 10, 1, 9, -39, -46, -71, -124, -149, -105, -30, -43, -76, -99, -7, 15, -29, -74, -17, -94, -89, -91, -78, -55, -99, -72, -48, 3, 11, 6, 35, 58, 61, 9, -49, -72, -98, -114, -84, -77, -55, -52, -11, 44, -18, -54, -101, -111, -111, -110, -89, -118, -124, -90, -30, -24, 16, 57, 77, 68, 62, 40, 25, -25, -30, -99, -86, -101, -83, -57, 35, 17, 9, -43, -65, -102, -96, -85, -61, -122, -96, -36, 11, 28, 44, 80, 111, 111, 109, 55, 52, 15, 28, -31, -59, -71, -66, -67, -13, 11, -6, -37, -109, -89, -106, -93, -28, 3, 2, 16, -4, 9, 52, 75, 111, 99, 60, 22, -1, 35, 61, 16, -36, -64, -69, -103, -52, 33, 12, -35, -45, 3, -18, 5, 43, 48, 89, 25, -18, -14, 34, 77, 94, 51, 12, -6, -31, 26, 23, 54, -12, -53, -59, -94, -55, -30, -11, -39, 47, 36, 51, 111, 27, 71, 75, 36, -7, -11, 2, 51, 31, 23, -59, -60, -20, 18, 27, 60, 31, -58, -30, -99, -70, -36, -6, 8, 98, 78, 115, 94, 70, 30, 33, -14, -25, -14, -19, 12, 38, -6, -71, -39, -20, 26, 39, 6, -42, -58, -48, -76, -101, -51, -15, 20, 43, 55, 46, 63, 39, 20, 26, 7, -14, -38, -14, -29, -1, -30, -37, -15, -3, 15, 10, -18, -62, -132, -60, -83, -105, -34, -14, -3, 83, 129, 73, 41, 23, 30, 11, -20, -35, 19, -42, -3, -1, -2, -18, -8, -9, 12, 25, -5, -53, -110, -117, -17, -25, -24, -15, 52, 48, 107, 81, 21, 2, -5, -40, 0, -5, -7, 0, 8, 30, 10, 20, 6, 27, 31, 3, -42, -42, -124, -90, -26, -38, -75, -14, -19, 36, 67, 37, -11, -32, -10, -18, -9, -3, -11, 0, 11, 5, 30, 65, 51, 58, -6, -28, -53, -90, -91, -69, -44, -21, -44, 9, -3, 23, 82, 23, 12, -33, -58, 9, 19, -7, -31, -35, 8, -6, 21, 36, 23, 10, -29, -46, -60, -95, -28, -61, -15, 16, 6, -16, -42, 7, 50, 8, -17, 10, 31, 24, -18, -32, -33, -57, -33, 8, 25, 45, -10, -31, -104, -108, -38, -22, -18, -44, -16, 16, -6, -20, -31, 37, 47, 49, 17, 35, 59, 29, 35, -7, 26, 11, -3, -8, -28, -42, -15, -29, -77, -72, -20, -25, -1, 38, 29, 7, 21, -13, 2, -30, -23, -24, 9, 37, -1, -33, 8, 40, -39, -32, -12, -23, -35, -51, -82, -95, -97, -76, 6, -40, -14, 15, -11, 43, -20, 12, -7, -16, -18, -49, -76, -55, -71, -28, 8, -17, -93, -105, -46, -45, -72, -25, -63, -79, -90, -28, 7, 0, -8, -3, -3, 8, 21, 13, 9, -6, -19, 11, -13, -30, -28, -26, -26, -4, -42, -42, -28, -2, 44, 15, 32, 13, 15, 6, 4, -18, -15, -8, -6, -11, -11, -15, -4, 8, -4, 11, -11, -2, -11, -17, 17, -2, 8, -12, 13, 3, 14, 13, -18, -19, -10, -15, -10, 13, 16, 14, -17, -1, -16, 12, -2647, -14, -9, 6, 0, 15, -42, -58, -52, -84, -82, -67, -15, 23, -23, -35, -47, -55, -54, -30, -6, -13, -16, -7, -10, -15, -4, 14, 1, -8, 9, -11, -16, -18, -4, 11, -40, -80, -59, -102, -40, 2, -61, -57, -88, -49, -33, -23, -61, -13, 6, 4, 30, 8, 19, -1, -8, -15, -7, 19, 6, 9, 3, -14, -55, -87, -97, -103, -86, -66, -93, -17, -26, -16, 2, 51, 73, 103, 69, 60, 2, -2, 29, -11, 11, -6, 23, 12, -67, -44, -48, -24, -65, -57, -30, 14, -12, -28, 11, -24, -15, -7, -7, 13, -8, 43, 24, -9, 58, 76, 1, 3, 12, 7, 51, -22, -56, -69, -74, -10, 0, 23, 48, 32, 22, 6, 6, -21, 9, -4, 24, -13, -53, -37, -45, 32, 57, 95, 35, -5, 9, 11, 11, -84, -99, -28, 10, 23, 27, 57, 17, 8, -9, -16, -8, -27, 0, -12, 2, -6, -9, 2, -35, 0, 37, 24, 14, 4, 11, -14, -41, -114, -73, -32, -2, -20, -2, 15, 0, -32, -20, 10, -4, 28, 31, 42, 80, 42, 80, 70, 48, 19, 44, 41, 17, -3, -15, 21, -44, -48, -19, -9, -10, 8, 44, 19, 20, 3, 15, -2, 5, 19, 45, 85, 78, 99, 110, 84, 73, 45, 30, 83, -2, 13, -5, -26, -60, -11, 12, -12, -16, 23, 21, 38, 31, -23, -8, 1, -30, -10, -28, 31, 58, 39, 47, 39, 60, 61, 86, 114, 23, -44, -13, -15, -40, -83, -5, -22, 26, 54, 44, 20, 0, -6, -4, -36, -81, -139, -176, -125, -87, -59, -52, -14, 27, 36, 81, 99, 22, 24, -39, -27, -49, -139, 14, 27, 1, 36, 26, 39, 36, -8, -11, -62, -145, -223, -325, -319, -291, -227, -144, -77, -50, 30, 67, 137, 20, 48, 10, -2, -54, -113, 57, 15, 32, 53, 44, 52, 39, 18, -26, -61, -40, -64, -115, -197, -210, -248, -212, -146, -73, -39, 66, 78, 8, 28, -16, -26, 28, -44, 53, 9, 28, 33, 28, 28, 6, 11, -7, -9, 25, 30, 36, -49, -80, -123, -134, -114, -71, -61, -15, 52, -10, 2, -4, -34, -19, -42, -11, -10, -16, 0, -14, -22, 14, -20, -17, 28, 31, 5, -3, -57, -49, -57, -22, -24, -38, -42, -4, 18, -76, -8, 2, -19, 7, -36, -78, -66, -65, 1, 12, 21, 40, 28, 8, -14, 51, 56, 14, 23, 13, 12, -9, -27, -24, 3, -35, -3, -107, -70, 17, 30, 46, -40, -185, -100, -79, -17, 9, 17, 61, 0, 1, 16, 51, 54, 67, 24, 23, -34, -54, -36, -52, -29, 11, -41, -75, -79, 4, 38, 40, 15, -121, -120, -81, -67, 9, -10, 39, 15, 8, -6, -2, 26, 19, -39, -60, -70, -79, -78, -45, -32, 38, 25, -61, -82, -3, 16, 45, 45, -82, -83, -33, -36, -48, -54, -39, -26, -17, -27, 8, -8, -25, -53, -44, -43, -39, -32, -23, -55, 8, 33, -20, -66, -20, 10, 55, 32, -84, -63, -18, -19, -73, -83, -57, -69, -50, -13, -9, -18, -31, -37, -27, -19, -15, 5, -15, -29, 31, -3, -46, -50, -14, 24, 24, -4, -97, -103, -15, -12, -29, -54, -26, -3, -16, -17, 4, -1, 9, -4, -21, -26, -20, -14, -52, -29, -9, -27, -50, -43, -4, 3, 32, 40, -62, -73, -24, -6, 30, -2, 28, 36, 26, -7, 15, 10, -10, -37, -7, -28, -26, -41, -15, 15, 8, -10, -52, 49, -11, 0, 82, 99, 5, -11, -44, -1, 21, 34, 48, 16, 37, -14, 13, -2, -24, -20, -8, -33, -8, -18, 0, 26, -4, -15, -21, 19, 12, -39, 70, 56, 30, 45, 13, -29, 35, 47, 12, 16, 22, 26, -6, 8, -35, -18, -29, -14, -14, 14, 28, 33, 10, 52, 13, -12, 17, -18, 64, 58, 23, -2, 2, -1, 2, 9, 42, -35, 8, 43, -12, 11, 8, 2, 14, 35, 44, 45, 33, 46, 14, 68, 22, 8, -5, 1, -21, -31, -4, -16, -27, 26, 39, -14, 7, -26, -29, 50, 17, 6, 53, 36, 50, 16, 31, 41, -7, 39, 47, 31, 40, 20, -18, 6, 10, -1, -33, -48, -92, -79, -27, 4, 2, 3, 50, 67, 48, 1, 12, 36, -9, -32, -75, -57, -37, -4, -6, -24, -11, -8, 20, 7, 18, -4, -3, 10, -1, -38, -55, -71, -58, -40, 6, 53, 8, -35, -35, -13, -18, -7, 0, -20, -3, 12, 19, 3, 0, 8, 2, -2, -7, -1, 12, 10, 17, 4, 15, 4, 0, -18, -5, -2, 1, 14, -16, -10, 11, 5, -14, -20, 5, 14, 12, -17, -1, -4, -8, 1216, -9, -3, -9, -17, -49, -24, -44, -27, -5, -28, -72, -33, 16, -7, -72, -2, 18, -22, -30, -23, 11, -8, 3, -23, -2, -10, 4, 16, -14, -17, 15, 20, 26, 1, 17, 45, 35, 23, 29, -18, -2, 52, 8, 5, 59, 31, -30, -27, -1, 12, 29, -1, -15, 19, 5, 15, -17, 5, -3, 78, 71, 57, 31, 43, 47, -7, 17, -31, 17, 11, 21, 19, -1, 33, 3, 29, 71, 50, 32, 1, -22, 23, -18, 2, 11, -29, -48, 35, 105, 73, 1, 35, 51, 27, -9, -7, 5, 20, 55, 37, 13, -16, -75, -39, 18, -3, -13, 34, 48, 2, 17, -20, 7, 37, 39, 35, 75, 68, 29, 57, 19, 10, 15, -11, -45, -2, 8, -24, -7, 26, 6, -10, -42, -50, 16, 72, 80, 30, -8, 15, 11, 10, 23, 40, 67, 15, 42, 32, 22, 7, 17, 0, -25, 9, -3, -33, -23, 0, -9, 16, -6, -15, -4, 39, 3, -36, 13, 10, 0, -56, 21, 2, -25, -14, 10, -17, -1, -14, 15, 4, 19, 16, 1, -9, -13, 0, 51, 41, 22, 25, 5, 20, -11, -20, -24, 0, 0, -82, 6, 20, 22, 14, -7, 12, -26, -13, -1, -18, -38, -32, 8, -28, -36, -21, 26, 5, -5, 30, 8, -7, 5, -28, 26, 19, -37, -84, -45, 29, 7, -23, -1, -20, -22, -23, -39, -74, -41, -14, -2, 35, 7, -5, -21, -9, -8, 11, 30, 18, 8, 2, -29, -2, -61, -71, -115, -4, -9, -23, -55, -17, -84, -105, -108, -94, -73, -4, 45, 81, 73, -5, -60, -20, -24, 48, 25, 9, 37, 34, -10, -27, -76, -109, -117, 1, 53, -30, -75, -65, -70, -117, -70, -58, -65, -14, 71, 74, 22, -49, -44, -31, -32, -8, 14, 53, 56, 10, 44, -9, -28, -102, -43, 7, 25, -50, -106, -79, -69, -95, -79, -69, -23, 51, 112, 59, 2, -12, -35, -65, -77, -56, 5, 55, 64, 23, 36, -15, -32, -51, 7, -5, -14, -76, -64, -51, -59, -35, -49, -18, 44, 97, 83, 70, 26, -3, -2, -44, -47, -42, -78, -2, 15, -47, 16, 11, -45, -57, 9, -22, -71, -57, -14, -27, -3, 9, -7, 30, 97, 153, 96, 54, -5, -22, -6, -21, -72, -55, -99, -45, -12, -66, 2, 14, -31, -12, 3, -24, -77, -48, 8, 15, 12, -9, -1, 57, 142, 154, 93, -5, -17, 9, 4, -3, -14, -63, -29, -2, 9, -87, -40, -4, -6, 53, 102, 8, -10, -26, 15, -6, 1, -27, 7, 89, 189, 96, -26, -54, -35, 4, 8, -29, 16, 15, 13, 51, -8, -105, -74, -22, 41, 102, 110, 114, 2, -18, -32, -23, -48, -53, 48, 122, 174, 70, -32, -37, 31, 9, 5, 21, 6, 41, 0, 8, -24, -116, -72, -44, 37, 85, 95, 101, 4, -30, -40, -52, -45, -51, -3, 66, 103, 25, -14, 19, 49, 33, 40, 38, 27, 23, -62, 2, -29, -98, -31, -27, 23, 81, 139, 88, 17, 7, 2, -14, -35, -26, 20, 56, 49, 17, 4, 11, 58, 17, 39, 46, 44, 22, -36, -27, -50, -19, -54, -20, 36, 49, 102, 75, 20, 32, -17, 0, -1, 8, 22, 44, 9, 6, -10, -5, 42, 18, -2, -1, -2, -36, -29, -51, -55, -90, -49, -22, 23, 28, 87, 48, 29, -11, -27, -8, 22, 0, 13, 22, 20, -5, -1, 24, 22, 24, -6, 9, -48, -54, -41, -55, -59, -81, 22, 16, 39, 92, 124, 89, 34, 25, -25, -1, -12, 10, 10, 39, 17, 49, 56, 64, 37, 11, 38, 20, -13, -43, -22, -24, -22, -44, 1, -5, 22, 80, 50, 15, 29, 14, 17, -5, -46, -52, -8, 3, 24, 46, 70, 47, 65, 24, 35, -15, -22, -9, -17, -34, 24, -22, 5, -18, -20, 84, 37, 49, -18, -13, 2, -34, -1, -17, -44, -19, 14, 44, 21, 6, 23, 15, -2, 1, -12, -29, -20, -27, 26, 14, 1, 6, -11, 3, 12, -17, -46, 5, 13, -3, -13, -7, -32, -22, 15, 3, -3, 29, -31, 9, 27, 24, -14, -21, 0, 41, 14, 6, 5, -4, 3, 16, -26, -34, -33, -23, -54, -24, 13, 31, 17, 47, 17, -51, -19, -38, -31, -72, -91, -27, -23, -21, 6, -6, 18, 8, 10, 6, -19, -2, -21, 5, -3, 1, -3, 16, -3, -12, -39, -25, -17, 16, -11, -10, -4, -9, 16, 4, -20, 14, 20, 8, -15, 3, 15, -13, 4, 13, 0, -15, 15, -2, -11, 11, 4, 7, -5, -12, -7, -16, -18, -3, -19, 20, 11, 1, 9, -20, 6, 2, -9, 3, -5, -20, -815, 10, 18, 10, 1, 2, 4, 19, 17, 16, 35, 61, 84, 57, 74, 66, 43, 30, 49, 59, 45, 35, 35, -5, 8, 19, 6, 4, 17, -17, 1, -9, 8, -24, 18, 16, 60, 59, 79, 52, 157, 144, 168, 85, 30, 42, 137, 138, 76, 96, 59, 50, 1, 6, 4, 15, -11, 4, -7, 24, 13, 8, 25, 9, 21, 11, -42, -29, -24, -23, -4, 13, 53, 33, 46, 92, 90, 93, 52, 135, 81, 13, -12, -1, -17, -6, -11, 1, -38, 12, -59, -19, -38, -86, -52, -22, -30, -32, -26, -23, -46, 19, 58, 8, 49, 77, 82, 121, 143, 69, 39, -6, -17, 10, 41, -16, -20, -40, -90, -84, -47, -55, -60, -47, -44, -19, 0, 2, 4, 46, 48, 4, 29, 69, 69, 96, 102, 50, 8, 6, -20, 8, -5, -60, -65, -63, -83, -55, -49, -22, -38, -50, -37, -35, -48, -8, 6, 25, 58, 32, 69, 40, 21, 35, 85, 60, 6, -12, 9, -8, -7, -7, -73, -58, -95, -60, -44, -29, -37, -56, -36, -40, -46, -17, -4, 24, 25, 19, 47, 26, 22, 30, 43, 60, 14, 0, 2, -12, 4, 31, -76, -81, -55, -36, -13, -19, -20, -33, -21, -47, -21, -65, -98, -43, -21, -16, -23, -3, -12, 7, 26, 90, -16, 12, 1, -15, 4, -2, -157, -77, -53, 9, -17, -23, -24, -13, -26, -54, -49, -117, -126, -143, -166, -154, -175, -126, -96, -38, 18, 75, 11, 38, -12, -22, 30, -13, -135, -69, -22, 33, -32, -22, -39, -33, -20, -38, -76, -120, -126, -172, -235, -305, -270, -222, -181, -118, -13, 40, 37, 20, 27, -6, 13, -26, -73, -31, 1, 33, 8, -30, -21, -28, -11, -2, -54, -27, -53, -78, -128, -199, -218, -202, -186, -141, -62, 29, 21, 41, 21, -22, -100, -151, -55, -53, 29, 46, 23, -10, 16, 26, -10, -11, 11, 17, 86, 52, 33, -24, -84, -107, -143, -86, -43, 17, 2, 57, -2, -35, 16, -134, -62, 31, 63, 78, 31, -13, 11, 25, 39, 43, 28, 44, 93, 105, 64, 32, -20, -59, -25, -40, -25, 18, 34, 43, -32, -43, -71, -82, -4, 10, 78, 65, 18, 16, 21, 34, 28, 38, 33, 56, 84, 45, 28, 39, 3, 22, -23, 1, -6, -4, 25, 15, -27, -35, -15, 28, 19, -27, 6, 37, -1, -3, 11, 32, 51, 49, 64, 59, 43, 39, 33, 14, -1, 29, 35, 20, 23, -24, 58, -20, -14, 35, 10, 46, -4, 41, 66, 26, 35, 7, 21, 40, 13, 36, 52, 37, 13, -7, 36, -17, -19, 49, -3, -22, 28, -23, 24, 6, 7, -22, 7, 52, -9, 61, 94, 53, 45, 19, 12, 57, 24, 12, 18, 4, -21, -7, -33, -68, 11, 14, 24, 15, 35, 73, 48, 29, 22, 1, 31, 84, -3, 22, 40, 58, 32, 10, -7, 11, 7, -26, -13, -32, -43, -18, -38, -10, 17, 14, 1, 15, 14, 75, 48, 33, 23, 17, 10, 40, -22, 3, 54, 27, 13, -6, 21, 23, -6, 26, 14, -33, 5, -6, 1, -11, 3, 27, 32, -18, 48, 25, 59, 71, 27, -26, -50, 14, -23, -41, 18, -4, -17, 1, 0, 18, 8, -3, -5, -3, 4, -4, -27, -2, 20, 11, 2, -10, 22, 24, 42, 51, -3, -11, 1, -11, -40, -68, -42, -34, -41, -11, -19, 16, -6, -36, 21, 4, 10, -26, 3, 14, -2, 10, 14, -14, 29, 58, 47, 72, -12, -6, -38, -77, -33, -88, -37, -42, -49, -24, -4, -19, 14, -23, -8, 14, -14, 25, 6, 14, 35, 3, 33, 20, 17, 49, 57, -11, 16, -19, -65, -56, -5, -15, -70, -61, -49, -37, 1, -38, -23, -17, -43, -3, -25, 3, -17, -7, 19, 41, 70, 65, 46, 23, -8, -11, -13, -15, -30, -7, -9, -64, -52, -49, -63, -3, 19, -68, -48, -16, -40, -33, -28, -37, -32, -55, -25, 5, 23, 28, 31, 28, 37, 8, 21, 20, -23, -26, 13, -34, -66, -31, -32, -38, 12, 9, -19, -16, 0, -16, 51, 24, -64, -40, -24, -26, 2, 20, -23, -4, 3, 6, 16, -11, -11, -15, -27, 10, 5, 0, 21, 5, -5, -18, -104, -91, -103, -129, -87, -43, -106, -85, -62, -74, -52, -27, 5, -8, -9, -4, -4, 9, -6, 8, 12, 0, -14, -15, -16, -24, -18, -22, -12, -23, -17, -41, -61, -30, -37, -28, -40, -60, -49, 3, -16, 9, -10, 20, 4, 1, -14, 14, 1, 16, 13, 12, -16, 18, -15, -12, -11, -1, -13, 4, 1, -3, -16, -4, -15, 6, -18, 4, 11, -7, -20, 6, -9, 262, 9, -18, -4, -18, 36, 19, 33, -8, 4, 29, 42, 22, 5, -31, -4, 6, 49, 52, 20, 63, 59, 54, 0, 2, 15, 14, 3, -8, -3, 16, 5, -2, 32, 75, 73, 26, 17, 31, 45, 105, 101, 52, 72, 71, 85, 51, 21, -20, 5, 37, 44, 12, -8, 19, -8, 12, 14, -7, 4, 41, 82, 96, 68, 1, 2, -18, 32, 19, 20, 13, 72, 76, 91, 70, 21, 51, 41, 80, 98, 80, 33, 9, -16, -4, -15, -8, -36, 10, 14, 7, 18, 0, -31, 5, 56, 57, 17, 10, -2, -51, -5, -34, -40, -24, -27, 6, 63, 82, 88, 26, 1, 7, 14, 42, -37, 15, -4, -6, 6, 5, 7, 18, 18, -2, -8, -8, -22, -51, -1, -40, -58, -101, -105, -49, -2, 6, 20, -3, 4, 19, 17, 25, -37, -25, 9, 14, -23, 3, 14, 4, -17, 8, -3, -18, -32, -45, -44, -25, -47, -89, -95, -127, -83, -42, -33, 0, 9, 9, 23, -63, -14, -28, -29, -24, -9, -31, -20, -7, -35, -12, -14, 0, -28, 2, -4, -5, -13, -12, -34, -73, -55, -42, -10, -14, 4, -7, 20, -36, 19, 16, -33, -31, -47, -45, -4, -11, 6, 21, 5, 19, 28, 23, 32, 56, 66, 58, -16, -17, 14, -31, 14, 12, 45, -7, -39, -78, -22, 41, -19, -40, -14, 23, 21, 20, -19, 16, -2, 8, 27, 67, 75, 92, 78, 104, 74, 37, 30, 11, 68, 48, 60, 8, -38, -30, -45, -34, -50, -14, 41, 13, 12, 23, 24, -2, -26, 1, -11, 15, 27, 80, 60, 74, 56, 31, 8, 0, 28, 44, -1, 38, -20, -27, -55, -11, -15, 38, 47, 37, 21, 10, -9, -35, -42, -56, -90, -80, -65, -45, -32, 0, 0, 36, 11, -16, 42, 31, 39, 10, -26, -71, -89, -34, 5, 34, 59, 45, 9, 39, -46, -100, -106, -149, -144, -123, -102, -119, -107, -18, 20, 43, 5, 11, -7, 37, 25, -2, -30, -48, -79, -35, 25, 64, 67, 55, -7, 10, -28, -77, -63, -122, -123, -73, -67, -85, -81, -28, 49, 70, 41, 18, -32, 17, 20, 28, -35, -46, -84, 4, 48, 59, 75, 29, 1, -37, -2, -27, -42, -94, -59, -24, -39, -40, -12, 33, 49, 29, 49, -3, -25, 20, 40, 1, -56, -31, -41, -46, -19, 21, 45, -16, -30, -22, -18, 3, -24, -14, -18, -14, 15, 21, 27, 71, 84, 48, 64, 35, -27, -15, -2, 11, -9, 41, -37, -47, -5, -22, -27, -16, -4, 47, 42, 36, 20, 17, 24, 58, 76, 64, 6, 60, 70, 1, -18, -14, 13, 21, 3, 3, 20, 21, 32, 38, 0, -32, -27, -21, -10, 29, 79, 76, 69, 41, 73, 54, 38, 21, -2, 9, -18, -27, -54, -25, -3, 58, -1, 33, -43, 24, 74, 78, 8, -19, -2, -13, -7, 13, -14, 18, 11, 7, 42, 19, 23, -5, 2, -20, -15, -47, -59, -44, 13, 5, 40, 30, 8, -4, 10, 29, -20, -34, -20, -10, -16, 7, -8, -14, -13, -9, -30, -26, -19, -40, -14, 7, -33, -54, -72, -24, -27, 4, 77, 23, -23, -10, 24, 48, 9, -32, -9, -19, -49, -22, -16, -11, -26, -14, -41, -38, -9, -38, -45, -31, -56, -58, 9, -66, -33, -22, 53, -23, 23, 14, 10, 29, 25, -8, -42, -18, -4, -10, -17, -6, -17, 29, -33, 0, 2, 8, -6, -33, -13, 17, 33, -24, -34, -28, 28, -11, -14, 42, 15, 66, 23, -9, -6, -21, -9, 3, -13, 19, -8, -14, -32, -29, -6, 4, -12, 4, 13, 15, 50, 30, 18, 7, 2, -5, -2, -1, -7, 15, 42, 10, -13, 6, 7, 14, -5, -21, -35, -26, -57, -49, -3, -19, 9, 7, 7, 42, 74, 37, -10, -16, -17, 17, -23, -3, 27, 56, 62, 49, 32, 34, 19, 21, 25, -29, 3, -21, -23, 6, 6, -4, 12, -13, -7, -4, 12, 71, 70, 12, 11, -5, 5, 10, 26, 0, -24, 7, 36, 62, 4, 17, 6, -7, 9, 11, 22, 38, 50, 38, 26, 31, 64, 22, 4, 24, 19, -2, -15, 16, -3, 6, -29, -35, -22, 54, 50, 59, 105, 50, 27, 42, 23, 32, 40, 50, 58, 10, 5, 4, 37, 35, 9, 41, 12, 20, -1, -19, -16, -10, -17, 19, 38, 60, 62, 78, 68, 34, 33, -9, 24, 0, 44, 85, 91, 71, 44, 22, 45, 36, 26, -6, -8, -3, -12, -19, -10, -16, -14, -19, -3, 16, -16, 15, 15, -5, 20, -7, 14, -15, -1, 5, 17, -12, -9, 9, -15, 16, -18, 8, 7, 10, 13, -13, 303, -19, 3, -14, 8, -12, -40, -12, -47, 20, 29, -24, 16, 35, 26, -15, 5, 27, -32, 5, -26, 12, 3, -14, -25, 8, -20, -10, 5, -6, 15, 4, 29, 33, -49, -11, -7, -43, 23, 58, 20, -12, 7, -9, 37, 46, -1, -17, 19, 57, 29, 23, 81, 32, -15, 3, 14, -3, -20, -2, 18, 3, -11, -7, 12, -11, 63, 47, 40, 7, -1, 7, -6, -7, -38, 2, -23, -6, -24, -37, -19, -19, 1, -16, 12, -3, -38, -16, -36, 0, -10, -60, -38, 23, 57, 28, 61, 27, -26, -32, -8, -41, -26, 17, -22, -37, -43, -55, -35, -53, -17, 18, 13, 6, -33, 20, -14, -8, -85, -72, -35, 4, 47, 11, 35, 19, -4, -39, -32, -47, -20, -23, 2, -48, -42, -1, -23, -30, -5, 17, -10, -11, -11, 7, -14, -54, -129, -96, -60, -24, 15, 21, 18, -6, -6, -8, -17, -18, -21, -21, -16, -30, -74, -23, -39, -33, -45, -14, 9, -13, -50, -32, -53, -73, -88, -102, -42, -1, 11, 10, -14, 0, 13, 20, -20, 4, -3, 47, -32, -45, -59, -89, -85, -79, -43, 12, 26, 23, -2, -40, -43, -56, -104, -75, -24, 5, 36, 23, 9, 33, 11, 26, 6, 15, 19, -15, -38, -79, -96, -124, -176, -128, -37, -20, -19, 7, -3, -54, -56, -48, -99, -68, -59, -19, -6, 4, -20, 4, 25, 46, 34, 47, 39, 10, -37, -79, -96, -125, -154, -82, -69, -19, 16, -1, -51, -82, -93, -81, -83, -79, -54, -75, -54, -14, -7, -9, 22, 58, 67, 51, 44, -9, -20, -82, -64, -128, -122, -43, -71, -13, -10, -43, -94, -64, -42, -43, -14, -51, -88, -90, -59, -25, -27, 35, 86, 36, 38, 34, 25, -14, -10, -29, -85, -80, -109, -41, -54, -15, -5, -46, -100, -22, -31, -19, -36, -86, -76, -78, -39, -22, 9, 33, 88, 42, 50, 6, -8, 3, 11, -23, -57, -101, -79, -28, 12, -10, -27, -36, -86, -16, -36, -28, 2, -57, -67, -7, 22, -8, 44, 26, 94, 41, 24, 16, 43, 19, 66, 14, -51, -74, -37, -13, 36, -18, 20, -44, -67, -28, 0, -14, 5, 11, 2, 0, 11, 27, 43, 47, 50, 44, -10, 25, 15, 28, 78, 22, -18, -84, -96, -67, -1, -7, 7, -39, -26, 6, 4, 59, 93, 89, 47, 60, -4, 12, 19, 48, 0, 11, -10, 33, 24, 63, 50, 66, -13, -83, -143, -110, -34, -24, 9, -18, -16, -8, 9, 80, 38, 60, 20, -6, 14, -2, -26, -56, -25, 23, 25, 57, 57, 58, 56, 18, 6, -92, -102, -112, -23, -8, -23, 3, 37, -3, -33, -23, -46, -18, -34, -28, -28, -53, -109, -104, -52, 2, 18, 42, 69, 77, 62, 15, -32, -89, -130, -89, -25, -34, -22, -30, -16, -42, -22, -14, -49, -42, -91, -59, -57, -90, -94, -80, -66, -19, -6, 15, 37, 29, 23, -32, -112, -164, -121, -74, -75, -25, -30, -44, 6, 33, -5, -22, -34, -25, -50, -53, -67, -31, -48, -23, -59, -10, -36, -25, -6, 27, 9, -15, -63, -126, -83, -76, -50, -26, -20, -3, 43, 54, 56, -10, -21, 4, -12, -21, -45, -31, -19, -24, -6, -15, -51, -21, -25, -27, -6, 5, -56, -40, -94, -80, -65, -70, -10, 26, 44, 79, 65, 48, 22, 55, 43, 7, 1, -35, -20, -2, -12, -32, -65, -45, -45, -1, 23, -33, -81, -47, -54, -60, -63, -25, -11, 48, 58, 121, 59, 48, 6, -3, 44, 24, 3, -16, -60, -31, -41, -83, -22, -33, -57, 5, 10, -1, -59, -50, -53, -37, -46, -3, 3, 52, 23, 43, 98, 34, -3, 5, 31, 21, -17, -28, -59, -81, -79, -83, -62, -68, -24, 4, 0, -55, -59, -42, -22, -22, 38, 2, -2, 27, 42, 7, 71, 106, 71, 26, 35, -8, 13, -14, -47, -47, -53, -71, -46, -62, 30, 66, 20, -17, -54, -34, -17, -16, -18, 11, -21, 9, 5, -13, 70, 123, 113, 74, 19, -20, 12, -16, -58, -9, -21, -19, -9, 17, 36, 41, 4, 55, 59, -13, -4, -8, -21, -9, -1, -2, 19, -29, -2, 58, 126, 65, 62, 68, 11, 43, 26, 54, 39, 42, 51, 59, 21, -21, 21, 69, 58, 37, 21, -8, 6, -4, -8, -17, -4, 1, 20, 6, 77, 65, 55, 43, 71, -3, -35, -7, 50, 40, 45, 57, 101, 56, 27, 62, 35, -5, 16, -8, -13, -3, -8, -5, -15, -1, -11, 11, 5, -11, -11, -13, -8, -11, -18, 11, -9, 20, 31, 2, -14, -15, 17, -7, -12, -10, 2, 20, -12, -16, -7, -647, -3, 13, 15, -15, 12, 16, 16, -4, 19, 42, 71, 28, 4, 38, 36, 0, 21, 44, 41, 50, 58, 53, -4, -10, 7, 2, -11, 17, 17, -3, -13, 8, 8, 49, 74, 85, 77, 83, 40, 44, 63, 90, 49, -9, 33, 129, 138, 77, 85, 33, -2, -49, 10, -9, 20, 20, 10, -21, -11, 21, 35, 33, 79, 65, 28, 2, 11, -13, 16, 81, 83, 139, 81, 99, 128, 148, 66, 44, 53, -6, 10, -17, 4, 18, -5, -38, -45, -2, 15, 0, 50, 36, 19, -16, 20, 4, -7, 17, 2, -11, 26, 54, 26, 51, 70, 99, 68, 84, 60, 20, 15, -2, -7, 44, -29, 33, -4, -9, -19, 9, 14, 8, 2, -26, -29, -34, 2, -7, 9, 23, -12, 20, 57, 69, 60, 80, 14, -14, -19, 19, 1, -7, -38, -30, -18, -36, -8, 3, -13, 6, -3, 4, -12, 17, -25, -21, -3, -3, -20, -6, 34, 57, 51, 32, -28, -23, 18, 9, -21, -50, -5, -11, -36, -42, -18, 27, 29, 18, -18, 10, -16, -20, -23, -16, -30, -51, -41, -18, 28, 45, 44, 6, -12, -42, -14, -20, -3, -5, 15, -3, 6, -2, -20, 22, 7, 1, 19, -8, -35, 3, -23, -42, -49, -57, -44, -4, 4, -4, 30, 36, -4, -62, -7, -13, -6, 23, 5, 9, 0, 5, -8, 6, 9, 0, 5, 15, -5, -6, -9, -63, -64, -38, -24, -21, -45, 13, 14, 4, 10, -11, 1, -3, 6, 52, -49, -57, 0, 49, 29, 32, 34, 31, 27, -23, -22, -5, -20, -50, -45, -33, -23, -5, -6, 11, -13, 2, -7, 38, 11, 28, -39, 16, -61, 22, 18, 4, 30, -24, 24, 11, 17, -7, -9, 1, -10, 4, -25, -28, 3, -15, 29, 4, -8, 13, 8, -17, 53, -1, 11, -29, -104, 13, 0, 22, -20, -32, -8, 25, -13, -44, -23, -34, 9, -48, -34, -1, 9, 0, -7, -12, -3, 39, 13, 0, 23, 19, -30, -32, -67, -3, 16, -27, -17, -17, -27, -8, -10, -15, 17, 16, 16, -67, -73, -30, -33, -42, -33, -15, -41, -13, -44, -15, 27, -9, -14, -7, -57, -4, -28, -68, -59, -32, -6, 15, 11, 22, 50, 39, 19, -57, -103, -61, -37, -37, -8, 11, -28, -13, 3, 16, -10, -20, -31, -21, -18, -11, -69, -48, -21, -2, -31, 2, 41, 66, 65, 99, 37, -38, -77, -60, -51, -41, 1, 8, -33, 45, 21, 25, -15, 18, 51, 67, 2, -84, -26, 7, -15, 18, 28, 27, 44, 70, 110, 122, 78, -3, -50, -42, -22, -17, -39, -52, 8, 37, 28, 15, -13, -11, 59, 74, 58, -50, 10, 30, 21, 53, 55, 43, 35, 63, 82, 124, 119, 36, 25, -22, -67, -6, -27, -9, -10, 65, 23, 20, -5, 7, 63, 84, 66, -58, -9, 50, 44, 66, 39, 26, 9, 8, 63, 118, 63, 35, 6, -11, -77, -45, -1, 31, 31, 12, 18, 22, 28, 1, 38, 67, 15, -55, 18, 52, 34, 21, -12, 14, 6, -32, 49, 87, 35, 34, -23, -2, -46, -3, 37, 13, 55, 70, 11, 21, 59, 30, 51, 34, -83, -54, -9, 36, 5, 12, 25, 9, -7, -21, 15, 74, 76, 29, -2, -22, -49, -7, 10, 40, 48, 51, 57, -16, 17, -14, -25, -6, -100, -63, -7, -6, 36, 57, 2, -17, 9, 6, 33, 49, 69, 33, 8, -8, -8, -31, -2, 16, 30, 62, 84, -21, 66, -12, -16, 19, -26, -61, -67, -12, 26, 48, -13, 26, -14, 14, 13, 47, 36, 41, 24, 8, -8, -8, 52, 77, 74, 16, 60, 1, -5, 3, -49, -2, -47, -42, -50, -5, 17, 15, 9, -1, 2, -29, -11, -13, 1, 2, -16, -16, 1, 10, 40, 27, 80, 29, 25, 0, 17, 5, -30, 2, -23, -5, -69, -23, 5, 8, 19, 18, -3, 10, 37, 15, -21, -34, -11, -14, -16, 2, -24, 32, 48, 0, 55, 20, 21, -4, -13, -3, -10, -8, -30, -55, -18, 37, 34, 9, 28, 34, 39, -14, 6, 24, -23, -3, -3, 23, 21, 2, 17, 7, 33, 41, 0, -7, -18, 5, 10, -2, -24, -49, -52, -20, 21, 8, 14, 25, 14, -34, -5, -2, -23, -48, -41, -73, -100, -82, -7, -29, -28, 4, -7, 5, -1, -20, -10, -11, -24, -59, -45, -74, -35, -81, -26, -12, -7, 36, -34, -41, -44, -44, -44, -47, -34, -27, 6, -19, -12, 14, 2, -8, -6, -12, 3, -16, 2, 7, 9, 1, -3, -12, -3, 20, 15, 18, -12, 4, -17, -11, -10, 8, -14, 4, 12, -11, -16, 7, 3, 14, -919, -19, -13, -19, -4, -26, 27, 50, 80, 87, 84, 92, 102, 75, 130, 93, 46, 37, 64, 46, 62, 30, 45, 13, 25, 9, -2, -5, -10, -13, 4, -16, 25, 8, 69, 69, 101, 120, 67, 65, 36, 43, 135, 98, 76, 68, 114, 91, 122, 118, 92, 73, 61, -15, 10, 13, -2, -15, 35, 35, -18, -35, 23, 15, 45, -8, -11, 26, 46, 18, 43, 30, 33, 24, 31, 70, 118, 67, 41, 79, 32, -20, -16, 7, 3, 1, 11, 85, 74, 29, 66, 0, -36, -77, -58, 0, -22, 24, -23, -3, -34, -36, -11, -27, 18, 42, 21, 9, -10, -78, 0, -20, 21, 0, -57, -23, 35, 32, 48, 7, -53, -83, -51, -6, -18, 17, 6, 1, 12, -17, -22, -45, -40, 7, 7, -24, -70, -69, -41, 15, 14, 20, -44, 14, 28, 23, 9, -3, -42, -61, -71, -53, 20, 46, 58, 40, 21, 26, 32, -24, -10, -23, 1, 33, -78, -40, -2, -21, -1, 21, 23, 46, 57, 8, 27, -13, -30, -44, -19, -6, 19, 61, 47, 44, 62, 58, 44, -4, 0, -5, 9, 56, 27, 21, 1, -6, 12, -8, 62, 95, 44, 32, -23, -43, -8, -19, -3, 8, 42, 60, 51, 44, 30, 41, 68, 19, 24, 44, 37, 35, 99, 56, 0, -24, -15, -3, 60, 52, 19, 13, 9, -7, -11, 14, 29, 13, 39, 24, 27, 21, 26, 64, 81, 62, 52, 70, 39, -14, 40, 24, 7, 43, 14, 15, 21, 52, 13, -1, 12, -19, -33, -1, 27, 13, 16, 45, -10, -53, -21, 20, 22, 38, 59, 108, 68, 19, 39, 52, -2, -17, 43, 75, 50, 38, -35, -48, -40, -31, -52, -5, 1, -2, 4, -20, -53, -68, -49, -33, -4, -17, 52, 30, 83, 78, 73, 41, -15, -5, 16, 52, 23, -9, -38, -66, -44, -17, -24, -29, -25, 10, -19, -37, -33, -25, -58, -54, -49, -31, -19, 5, 50, 93, 110, 25, -19, -30, -8, 35, 32, -28, -27, -93, -45, -17, 19, 17, -2, -12, -9, 21, -8, -8, -64, -73, -36, -49, -42, -10, 10, 54, 48, -7, -37, -29, -14, 32, 39, -54, -33, -12, -16, 0, -7, 11, 5, -30, -1, 36, 28, -4, -39, -66, -25, -41, -48, -12, -24, -16, 48, 47, 6, 0, -7, 53, 42, -16, 8, 17, -19, -43, -28, 7, 12, 27, 17, 1, 55, 1, -102, -60, -43, -35, -64, -31, -43, 10, 85, 39, 50, 5, -8, 44, -17, 13, 27, 46, 34, -2, 16, 23, 67, 49, 14, 3, 68, -33, -105, -111, -100, -55, -28, -65, -36, 30, 46, 35, 49, 22, -10, -6, -101, -34, 35, 79, 73, 74, 49, 29, 77, 58, 31, 36, 97, 31, -60, -100, -93, -62, -28, -36, -25, -3, -13, 40, 41, 49, 4, 22, -51, -75, -30, 29, 39, 12, 15, 50, 44, 57, 49, 57, 192, 115, -42, -61, -77, -49, -25, -47, 4, 34, 1, 50, 54, 18, 20, 33, -30, -121, -45, -33, -3, -2, 10, 33, 26, 22, 10, 78, 137, 100, -6, -30, 3, -62, -55, -46, -51, 14, 3, 51, 25, 27, -8, -34, -82, -145, -119, -39, -6, -1, 29, 6, 18, 22, -1, 59, 98, 42, 11, 9, -51, -74, -57, -54, -25, -29, 11, -22, 6, 33, 11, 25, -65, -63, -94, -31, 5, 41, 61, 32, 24, 16, 27, 57, 91, 33, 35, -12, -31, -56, -72, -50, -48, -28, 3, 31, 20, 22, 21, -8, -57, -58, -72, -56, -24, 66, 59, 41, 64, 36, 77, 58, 63, 50, 10, -2, -11, -27, -68, -63, -35, -28, 6, 24, -18, -4, 6, -18, -8, -51, -16, -49, -67, 12, 26, 32, 39, 0, 37, 30, 39, 37, -9, 26, 3, -41, -36, -70, -24, -11, 24, 8, 26, 17, 12, 0, -28, -38, -63, -62, -48, -57, 1, 11, 37, 55, 43, 25, 42, 51, 13, 17, -2, -35, 2, -3, 9, -27, -13, 2, -10, -6, 9, -9, -2, 19, 25, 6, -68, -42, -9, 31, 76, 112, 107, 53, 59, 65, 40, 4, 3, -5, -16, -33, -12, -2, -25, 46, -3, 19, 8, -8, 14, 41, 36, 25, -7, 10, 5, -26, 2, 25, -9, -28, -43, -31, -33, -18, 21, 7, -15, -26, -17, -18, 24, 38, 9, 9, 17, 13, -2, -16, -5, 39, 35, -7, 17, 9, 13, 12, 69, 15, -16, -26, -5, 22, -29, -19, -26, 7, 38, -5, -9, 0, -2, 2, -17, -8, -6, -1, 12, -20, -15, 18, 10, 17, 13, 12, 1, -8, -9, -8, 3, -13, -7, 11, 10, -20, 11, -6, 10, 19, 4, 1, -7, -1643, 3, 18, -12, 18, 41, 52, 44, 45, 46, -16, 12, 23, -25, -27, 2, -8, -15, 21, 33, 16, 7, 15, 21, -1, -18, 1, 2, 9, 11, -20, 20, 11, -11, 39, 6, -14, 29, -26, -58, 11, 8, -41, 26, -13, -41, -8, -58, -26, -37, -60, -51, -53, 11, 12, -13, 19, -11, -16, -4, -3, -72, -48, -70, -94, -57, -118, -121, -82, -85, -59, -43, -58, -48, -71, -60, -42, -61, -48, 11, 21, 18, 6, 3, 13, 7, 37, -6, -25, -125, -119, -79, -131, -95, -44, 3, -38, 41, 42, 53, 30, -7, 0, 5, -16, -31, -17, 15, 8, 21, 12, -7, 17, 5, 67, -20, -29, -116, -98, -90, -93, -59, -36, 5, -4, 43, 49, 58, 95, 78, 42, 43, -1, 8, -18, -30, -93, -66, -12, -10, 20, -6, 51, -19, -49, -32, -38, -57, -68, -10, -20, 6, 47, 74, 50, 64, 74, 34, 62, 30, 29, 6, 7, -24, -87, -60, -55, 0, 9, -12, 26, -3, 26, -28, -55, -55, -7, -18, -3, -11, 25, 39, 62, 40, 48, 48, 37, 33, -12, 27, -28, -41, -55, -21, -15, -28, -7, 20, -21, 5, 6, -51, -59, -42, -25, -22, -38, -18, -27, -8, 36, 77, 113, 94, 62, 24, 10, -4, -26, -41, 8, -23, 39, 44, -4, 22, -32, 14, -24, -21, -9, -21, 8, -16, -17, -4, -34, 5, 33, 47, 85, 43, 28, 12, 2, -24, -46, -45, -14, -74, 46, 64, 12, -12, 13, -7, -24, 6, 36, -2, -2, 9, -29, -4, -17, -22, -11, 4, -7, -35, -35, -24, 14, -22, -67, -29, -27, -84, -49, -7, 23, 38, -15, 17, 16, 29, -4, -26, 16, 15, -36, -41, -27, -45, -27, -32, -76, -61, -40, -45, -23, -27, -69, -40, -4, -88, -25, 26, -20, -6, -57, -17, 50, 24, 9, 14, 51, 11, -38, -77, -73, -57, -70, -69, -94, -54, -69, -20, 14, 9, -51, -37, 18, -72, 8, 9, 15, -63, -84, 39, 87, 55, 3, 45, 44, -19, -48, -67, -90, -72, -100, -84, -37, -58, -60, 2, -10, 22, -44, 1, -32, -55, 42, -1, -9, -45, -74, 24, 72, 62, 30, 55, 31, -5, -31, -86, -106, -91, -108, -94, -43, -11, -10, 23, 41, 8, -13, 1, 2, 2, 69, -10, 31, -55, -78, -13, 48, 56, 33, 28, 6, 14, 22, -49, -99, -95, -60, -40, 15, 23, 72, 41, 55, 27, 38, 35, 31, 17, 61, 2, 7, 46, -29, 13, 7, 34, 27, 25, 24, 49, 42, 18, 7, -21, 2, 32, 54, 66, 47, 55, 48, 59, 10, -24, 7, 47, 67, 43, 10, 23, -67, -24, 19, 11, 62, 56, 60, 36, 69, 66, 31, 51, 70, 84, 37, 37, -3, -9, 10, 32, -2, -20, 14, 54, 81, 61, 31, -39, -35, -13, 33, 6, 22, 42, 19, 0, 32, 88, 89, 80, 56, 79, -8, -42, -14, -8, -11, -18, -4, 20, -9, 22, 46, 40, 16, -8, -67, -40, 7, -16, -23, -30, -39, -33, -6, 26, 79, 64, 32, -11, -69, -69, -24, -11, 3, 10, 2, 9, 59, 11, -20, -2, -4, -23, -63, -72, -57, -35, -27, -11, -13, -57, -32, 42, 30, 3, 14, -40, -56, -77, -31, -5, 1, 8, -23, -5, 50, 47, -9, 47, 16, 2, -54, -92, -53, -17, -25, -33, -23, -16, 16, 15, -23, -34, -10, -15, -27, -3, 18, 8, -31, 12, 31, 12, 54, 58, 2, 18, 2, 31, -65, -122, -65, -26, -6, 2, -7, -19, 20, -7, -11, -17, 16, 29, -17, 15, 18, -7, -14, 17, 69, 72, 51, 54, -24, -16, 1, -32, -41, -116, -95, -20, -20, 0, 12, 13, 47, 11, 43, 43, 18, 34, -18, -4, 30, -4, 4, 23, 40, 45, 31, 5, 34, 5, 2, -30, -74, -97, -123, -30, -14, -6, 8, 32, 23, -8, -14, 32, -4, -23, -46, -37, -66, -46, -17, 13, 13, 50, 44, 48, 38, 3, -1, -10, -11, -55, -34, -35, -45, -26, 52, 40, -15, 16, 14, 19, -14, 2, -22, -21, 14, -3, 79, 48, 51, 7, -19, 48, 22, 16, 16, 5, -18, 32, 65, 102, 73, 86, 87, 60, 35, 22, 72, 109, 34, -3, -12, 31, 14, -14, 51, 60, 62, 37, 29, 43, -12, 15, 5, 21, -2, 6, 10, 30, 66, 66, 57, 52, 118, 41, 26, 64, 11, 53, 78, 61, 26, 42, 27, 52, 24, 19, -14, 19, -4, 16, -15, -18, 12, -15, 16, -3, -4, -6, 16, -18, 2, 6, -16, -2, 7, 14, -6, 5, -1, 6, 5, 16, -1, -1, -2, 20, 12, -6, 1, -1503, -6, -6, -7, -11, 29, 44, 54, 63, 66, 68, 74, 101, 88, 122, 81, 25, 28, 39, 67, 60, 24, 20, 24, 22, -2, 4, 3, -12, 16, 19, 2, 22, 33, 66, 80, 116, 112, 107, 111, 94, 76, 171, 118, 78, 105, 110, 121, 93, 118, 78, 54, 70, -4, 19, -5, -1, 2, -5, 13, -31, -37, 11, 61, 64, 54, 34, 36, 44, 9, 37, 48, 32, 21, 35, 61, 69, 65, 41, 90, 29, -36, 30, 6, 4, 12, -38, -61, -3, -12, -11, -5, -22, -16, -18, 44, 25, 55, 11, 42, 36, 37, 67, 45, 74, 80, 42, 27, 92, 47, 29, 14, 2, -11, -24, -76, -21, -20, -20, -49, -79, -54, -14, 33, 29, 53, 32, 49, 37, 59, 49, 19, 52, 48, 27, 26, -27, 32, 3, 20, 3, -15, -11, -62, -45, -55, -61, -75, -77, -88, -18, 17, -5, 20, 51, 13, 7, 10, -12, -2, 38, 46, 79, 27, -30, -19, 4, -19, -10, 22, -11, 4, -24, -110, -78, -48, -71, -41, -23, -21, 21, -2, -35, -14, -10, -3, 20, -12, 15, 40, 76, 63, 6, 34, 15, 23, -21, 16, -32, 41, 26, -34, -74, -69, -54, 8, -17, -20, -32, -1, -12, -19, -6, -32, 5, 24, 34, -2, 4, 28, 42, -12, -27, 25, -12, -29, -22, -14, 24, 1, -9, -47, -37, 11, -16, -13, -39, -48, -53, -14, -2, 11, 41, 9, 3, -3, -51, -38, -17, -17, 11, 49, -9, -15, 16, 19, -26, -8, 23, -39, -48, 3, -21, -27, -49, -13, -40, -54, -11, 45, 58, 37, -2, -32, -36, -22, -37, -2, 13, 3, 49, 53, 7, -19, 54, -20, 16, -46, -66, -15, -38, -50, -61, -56, -55, -30, 7, 42, 26, 39, -18, 0, -17, -30, -35, -14, -28, 39, 7, 6, -65, -57, 28, 9, 2, -49, -15, -7, -11, -56, -72, -86, -87, -51, -8, -3, 15, -19, -21, -46, -19, -17, 20, -37, -31, 23, 12, -12, -35, 9, 56, 18, -3, 12, 44, 24, -27, -65, -79, -45, -60, -16, -49, -26, -47, -36, -53, -44, -15, 5, -18, -37, -66, 18, -8, -19, -33, 38, 17, 2, 19, 68, 64, 20, -2, -43, -41, -57, -32, -35, -52, -50, -30, -63, -41, -48, -43, -27, 19, 35, 47, 26, -26, -11, -4, 38, 7, 3, 20, 38, 26, 30, -12, -10, -46, -42, -21, -55, -64, -52, -60, -50, -40, -34, -54, -31, 47, 50, 28, -12, 2, 43, 23, 30, 6, 62, 67, 45, 46, 47, 26, 33, 22, -2, 32, 4, -45, -36, -21, -42, -30, -27, -14, -16, 50, 37, 39, 16, 22, 61, 22, 28, 9, 48, 87, 27, 61, 31, 44, 36, 20, 71, 93, 91, 48, 15, 2, -9, 32, 16, 20, -20, -2, 22, 59, 16, -13, 61, -8, -19, -37, 7, 40, 4, 6, 9, 35, 35, 34, 25, 119, 96, 16, 14, 9, 18, 5, 11, 27, -18, -43, 21, 55, 10, 14, 41, -37, -39, -8, 12, 10, -25, -29, 43, 37, 31, 31, 86, 80, 67, 33, -7, 28, 10, 7, 0, 14, -9, -6, 28, 32, 63, 7, -7, -14, -67, -54, -13, 34, 15, 7, 64, 62, 67, 63, 85, 75, 59, 50, 13, 0, -4, -14, 7, 3, -39, -4, 27, -12, 11, 17, -22, -58, -33, -9, 8, 16, 28, 64, 73, 69, 86, 72, 72, 93, 65, 20, -30, -7, -10, -27, 5, -24, -35, 1, 33, 6, 12, -16, -21, -32, -48, -40, -35, 41, 74, 87, 74, 103, 83, 64, 48, 61, 59, 3, 14, -18, -20, -13, -5, -5, -13, -7, 45, 13, -11, -1, -54, -16, -8, -48, -3, 8, 33, 32, 34, 17, 30, -23, 17, -21, 21, -27, -17, -58, -51, -42, -13, -2, -8, -34, -11, 5, 14, 14, -21, 29, -8, -26, -57, -4, -33, 23, 20, -7, -20, -36, -10, -21, -22, -24, 13, -51, -44, -37, -51, -57, -51, 0, 36, 15, 6, 0, 17, -20, 14, -31, -45, -54, -38, 23, -14, 8, 31, -2, -16, -4, -30, 26, 12, -46, -67, -31, -7, -38, -16, -40, 26, 8, -19, 10, -10, 15, 16, 11, -26, -58, -94, -70, -33, -40, -33, 10, -26, -35, -1, -32, -22, -41, -48, -21, -13, -21, -17, 14, 15, -11, -18, 2, -1, 18, 9, -18, -6, -29, -21, -37, -10, -45, 29, 48, 67, 35, 37, 20, 24, 3, 5, -31, -10, -3, -7, 12, 2, -13, -20, 5, -13, -13, -11, 19, 0, -3, 0, 3, -16, 7, 16, 4, 14, 5, -21, 9, 11, 2, 10, 12, 3, 16, -18, 0, 9, -2, -18, 9, -1500, 16, 12, -14, -15, 17, -34, -18, -43, -28, 10, 24, 35, 4, -61, -4, -10, -15, 7, -14, -11, -36, -18, 14, -14, 5, 7, -4, 0, 14, -4, 20, 3, -19, -62, -95, -133, -91, -82, -64, -44, -17, -73, -70, -57, -41, -69, -38, -30, -50, -55, -34, -49, -24, -7, -14, 12, 6, 2, 22, -69, -15, -141, -134, -140, -98, -58, 0, 39, -32, -6, 9, 10, 19, 5, 34, 38, 33, 6, 32, 41, -31, -35, 9, 3, -7, 13, 37, -24, -46, -60, -72, -53, -84, -14, -17, -4, -27, 29, 33, -9, -10, -11, 6, 24, -15, -12, -36, 37, 41, 63, -19, -15, -2, -5, -7, -51, -38, -57, -23, -26, -9, 5, -10, -3, -21, 6, 24, -46, -56, -36, -28, -36, 28, 30, 15, -16, 16, 75, 12, 14, -7, -21, -24, -23, 7, 8, 20, 0, 39, -16, 12, -14, 0, -3, -16, -30, -4, -36, -13, 8, 18, 2, 12, -7, 42, 100, -13, -11, -5, -10, -31, 4, 12, -19, -7, -10, 15, -2, -11, -12, -8, -30, -24, -52, -39, -33, -5, 20, 14, 5, 11, 32, 109, 88, 10, 9, -31, 46, -25, 1, -27, -43, 14, 11, -31, -10, 4, 10, -11, -6, -10, -78, -41, -33, -11, -10, 15, 37, 39, 67, 83, 22, -27, -19, 14, 48, 45, -20, -58, -29, 17, -29, -31, -43, -4, 16, 17, 4, -19, -89, -50, -51, 2, -15, 30, 27, 67, 52, 70, -19, -29, 16, 0, 50, 36, -11, 19, 3, 6, -11, 3, -4, 19, 14, 16, -7, -18, -3, -23, -54, -10, -1, 24, -4, 46, 36, 69, 91, 31, -43, -1, 79, 34, 7, 21, 17, 36, -1, 52, 49, 17, -11, 7, -10, -19, 3, 3, -10, 5, 2, 48, 24, 57, 70, 58, 63, 48, -13, -14, 110, 42, 40, 45, 15, 93, 45, 77, 54, 17, 16, 29, 33, 43, 46, 16, -4, 37, 51, 45, 51, 42, 72, 37, 64, 28, -3, 28, 113, 1, 16, 54, 53, 70, 3, 36, 40, 18, 22, 9, 8, 25, 33, 12, 17, 14, 14, -15, 38, 57, 40, 23, 86, 12, -25, 24, 80, 90, -18, -29, -16, 24, -20, 7, -6, 34, -15, -30, 12, 13, 27, 46, 6, 1, -46, -36, -47, -37, 10, -43, 74, 34, -8, 28, 98, 85, 55, -59, -37, -6, -59, -65, 10, 21, 12, -24, -51, -20, 13, -9, -34, -50, -51, -113, -87, -121, -113, -56, 61, 42, 15, 11, 46, 67, 30, -77, -64, -72, -66, -43, 2, 37, 34, -19, -60, -37, -6, -72, -71, -120, -103, -117, -140, -110, -89, -11, 45, 20, 8, -29, -4, -5, -88, -165, -151, -101, -43, 16, 39, 90, 60, -18, -102, -133, -91, -90, -81, -107, -109, -83, -101, -53, -31, 45, 50, 22, 20, 21, -24, -86, -214, -167, -117, -63, 13, 68, 100, 88, 34, -89, -180, -125, -78, -37, -26, -58, -17, -57, -42, 13, 22, 80, 89, 40, 13, -29, -55, -132, -198, -107, -38, 15, 16, 48, 83, 96, 13, -117, -168, -65, 35, 36, 34, 34, 12, 10, -22, 45, 28, 63, 78, 35, -1, 5, -58, -176, -211, -87, 1, 7, 42, 102, 97, 75, -3, -84, -64, -13, 71, 74, 47, 14, 2, 21, 46, 35, 65, 61, 48, 32, -25, 20, -50, -179, -132, -46, 16, 76, 92, 134, 83, 23, -46, -125, -78, -2, -5, 20, 30, -1, 18, 30, 60, 46, 96, 90, 11, 87, 15, -9, -15, -100, -62, -12, 1, 68, 91, 73, 35, 5, -56, -147, -132, -67, -42, -13, 12, 52, -13, -2, 16, 50, 36, 69, -10, 23, 20, -54, -70, -40, -66, -6, 30, 24, 49, 30, 16, -34, -39, -85, -108, -72, -16, -16, -1, -11, -15, 1, -15, 2, 5, 24, 10, 14, 7, -37, -81, -89, -80, -137, -44, -36, 6, 41, 35, 23, 43, -16, -18, -11, -4, -1, 0, -46, -63, -5, -36, 21, -40, -15, 20, 1, -19, 17, -30, -42, -73, -94, -63, -28, 4, 28, 27, 42, 73, 45, -16, -70, -57, -48, -72, -66, -99, -98, -30, -24, -57, -49, 0, -18, 9, 6, -20, 25, -26, -63, -75, -30, -21, -28, -13, 16, 64, -7, -27, -29, -87, -117, -109, -82, -76, -71, -27, -37, -60, -17, -17, -10, -9, 13, 10, 1, -12, -28, -59, -49, -64, -40, -75, -52, -17, -21, -18, -80, -91, -76, -67, -27, -27, -54, -39, -27, 14, 16, -13, 0, -9, 5, 9, 8, 10, 12, 0, -9, 15, -8, -1, 7, -5, 17, -8, -25, -10, -13, 3, -2, -14, 6, 12, 3, -17, 0, -16, 9, 1, -1781, -8, -6, 0, -17, -23, -43, -52, -39, -3, -11, -26, -56, -49, -81, -61, -60, -53, -59, -50, -24, -28, -41, -13, -7, -14, -5, -18, 19, -20, -3, 5, -34, -18, -13, -41, -49, -28, -91, -96, -73, -103, -131, -108, -149, -84, -130, -121, -99, -85, -12, 13, 9, -19, -6, -1, 5, 6, 11, 13, -40, -47, -77, -88, -71, -86, -129, -162, -191, -167, -146, -134, -130, -94, -107, -112, -121, -76, -62, -31, -23, -25, 0, 1, -12, -9, 16, 42, -20, -57, -64, -10, -31, -79, -65, -35, -21, -10, 0, 8, -14, -17, -48, 27, 11, -25, -18, -12, 6, -18, -6, 3, 11, 10, -7, -39, -47, -71, -61, -34, -35, -20, -9, 26, 39, 39, 13, -5, 23, 0, 13, -7, 4, -12, 15, -9, 11, 5, 31, -11, -10, -1, -14, -36, -52, -22, -42, -18, -42, 18, 10, -4, 39, 26, 3, 33, 23, 3, 20, 6, -5, -27, -16, -12, -4, 38, 66, 23, -3, -7, 31, -12, -23, 3, 9, -16, 18, 37, 35, 8, 11, 20, 39, 26, 33, 37, 60, 40, 18, -7, -18, -13, 9, 48, 1, 8, 4, 6, 41, -18, -29, -25, -3, 37, 24, 46, 43, 11, 14, 31, 43, 52, 61, 72, 55, 71, 14, 46, -14, 28, 46, 49, 8, 24, -1, 38, 8, -17, -27, -2, 26, 16, 51, 30, 24, 23, 13, 34, 74, 42, 79, 61, 73, 75, 40, 46, 27, 33, 65, 57, 3, -3, 9, 46, -46, 89, 33, 2, 51, 49, 1, 60, 78, 13, 32, 32, -1, 17, 34, 39, 65, 91, 92, 77, 28, 56, 93, 95, 6, -16, -19, 39, 26, 64, -14, -5, 48, 41, 50, 87, 66, 16, 8, -26, -17, -32, -12, 35, 39, 67, 69, 69, 56, 101, 63, 58, 2, -34, 16, 54, 88, 58, 43, 44, 40, 73, 100, 107, 39, -24, -51, -43, -58, -48, -24, 16, 12, 3, 37, 45, 68, 103, 99, 38, 21, -20, -19, 7, 19, 41, 52, 31, 14, 35, 66, 38, -7, -32, -67, -76, -78, -59, -51, -34, -39, -26, 16, 47, 67, 70, 46, -11, 26, -5, -22, -10, 4, 18, 49, 57, 21, 40, 7, -5, -17, -67, -50, -64, -72, -82, -50, -45, -44, -17, -5, 9, -4, 17, -14, -24, -40, -8, 5, 4, -55, -15, 42, 36, -12, 1, -33, -32, -3, -41, -13, -23, -40, -40, -56, -76, -56, -57, -39, -30, 1, -35, -54, -18, -58, 2, -12, -57, -96, -62, 37, -19, -30, -13, -33, -38, -17, -13, 0, -3, 11, 9, 12, -48, -53, -42, -70, -89, -62, -65, -75, -25, -29, -7, -7, -22, -143, -116, -24, -2, -53, -27, -10, 25, -23, -3, 30, 27, 50, 29, -6, -67, -65, -103, -85, -85, -74, -77, -66, -24, -14, 10, -14, -41, -119, -146, -57, -47, -61, -30, -27, -44, -22, 15, 44, 70, 63, 36, -17, -26, -79, -57, -96, -65, -72, -32, -29, -36, 3, -35, -9, -75, -122, -144, -70, -77, -69, -12, -24, -35, -37, -22, 9, 42, 22, 36, -15, -52, -47, -63, -88, -80, -54, -15, 15, -31, -15, -35, -12, -38, -40, -200, -124, -87, -53, -16, -19, -19, -65, 6, 31, 21, 42, 21, 23, -13, -63, -53, -91, -55, -43, -42, 17, -31, -34, -20, 32, 12, -23, -85, -43, -59, -20, -25, -1, -20, -41, -19, -8, 19, 45, 46, -18, -4, -41, -68, -66, -19, -15, -3, 36, -4, -14, -15, 15, 21, -40, -58, -23, -30, -21, -3, -28, -51, -24, 13, 22, 31, 14, 22, 6, -30, -30, -36, -52, -25, -3, 23, 58, 16, -1, 5, 14, 21, 10, -16, -23, -39, -52, -43, 5, 3, 2, 28, 20, 41, 43, 27, -10, 9, 27, 22, 38, -2, 5, 6, 61, -18, -29, 9, -9, 10, -19, -41, -39, -28, -50, -37, -8, -28, -33, 15, 34, 46, 49, 36, 62, 50, 93, 130, 84, 36, 31, 11, 2, -25, -8, -14, 12, 17, 23, 24, 14, -12, -45, -9, -6, -23, -19, 39, 57, 64, 127, 133, 140, 193, 159, 169, 118, 116, 85, 49, 36, 39, -39, 14, -6, -8, -3, -8, 16, 77, 44, 78, 13, -5, -26, 40, 64, 103, 151, 162, 181, 128, 91, 114, 97, 80, 52, 36, 17, 5, 5, 4, -20, -5, -9, -20, 20, 35, 42, 42, 71, 41, 69, 59, 50, 10, -29, 79, 79, 56, 62, 26, 42, 54, 33, 2, -10, 18, 11, -6, 1, -11, 17, -3, -11, 19, 11, -14, 11, 0, 13, 15, -1, 13, 16, 19, -3, -3, 16, 20, -18, 1, -5, 14, 8, -20, -12, 7, 7, -1185, 3, -7, -8, 20, 14, 64, 72, 49, 57, 41, 104, 144, 114, 127, 43, 3, -2, 30, 77, 59, 32, 51, 20, -4, 3, 7, -20, -18, 0, 8, 9, 1, -25, 28, -2, -5, 6, -13, -12, 23, 29, 96, 35, -23, -19, 38, 46, 27, 54, 58, 21, 50, -7, 9, 10, -5, -6, -23, 3, -47, -7, -10, -23, -46, -49, -48, -72, -51, -32, -19, -57, -34, -27, -36, -4, 17, 4, -13, 47, 31, 37, 0, -2, -2, -15, -24, -32, -64, 18, -14, -19, -26, -66, -64, -77, -61, -46, -58, -25, -31, -21, 13, 4, 10, 46, 24, 51, 14, -27, -12, 1, 16, -13, -17, 2, -3, -7, -25, -7, -54, -18, -41, -43, -39, -39, -34, -22, -30, -12, 2, -11, 27, 79, 54, 10, -15, -86, -86, -18, -12, 13, -39, -5, -20, -33, -16, -26, -76, -49, -63, -28, -52, -28, -32, -37, -28, -7, 20, 34, 38, 53, 57, 39, -30, -80, -67, 4, 9, -16, -56, -5, 7, -40, -36, -58, -111, -81, -61, -71, -39, -38, -78, -43, -66, -37, -2, -9, 13, -40, -37, 18, -51, -94, -54, 6, -13, 13, -44, -7, -35, -70, -49, -82, -128, -80, -75, -49, -37, -60, -59, -74, -69, -75, -66, -67, -88, -88, -52, -41, -60, -70, -17, -9, -10, 26, -40, -10, -123, -163, -140, -113, -116, -91, -93, -56, -44, -22, -17, -65, -77, -59, -78, -83, -66, -49, -83, -65, -88, -36, 4, 5, -1, -18, 18, -60, -124, -141, -128, -75, -69, -68, -48, -22, -7, 21, -4, -19, -38, -47, -35, -51, -35, -54, -88, -97, -74, -86, 1, -7, 4, -84, -47, -57, -57, -87, -41, -46, -43, -24, 14, 26, 28, 34, 31, 33, 2, 3, 15, 29, 37, -23, -52, -63, -63, -65, -10, 4, -16, -55, -95, -139, -125, -74, -42, -15, -32, 37, 31, 64, 35, 56, 53, 0, -8, -27, 6, 15, 72, 10, -15, -33, 3, -7, -37, 26, -3, -25, -59, -119, -142, -30, -25, -25, 9, 56, 65, 84, 39, 78, 11, -9, -41, -17, 25, 9, 37, 12, -40, -35, 10, 59, 5, 11, -2, -22, -104, -47, -66, -74, -56, -50, 35, 89, 83, 76, 48, 52, 19, -21, -31, -39, -10, 11, 28, 21, -32, -24, 79, 76, 64, 44, -24, -54, -43, -20, -95, -106, -47, 10, 18, 62, 41, 33, 82, 80, 22, -60, -71, -17, 4, 26, 34, 30, -10, -58, 25, 68, 69, 10, -13, -5, -27, -39, -67, -84, -62, -5, 7, 43, 70, 71, 84, 82, -15, -60, -23, 30, 14, 9, 60, -1, -34, -85, -29, 25, 67, 18, 26, -1, -65, -74, -107, -113, -29, -15, 31, 23, 36, 70, 69, 74, -32, -76, 23, 34, 31, 6, 24, -28, -18, -55, -30, 18, 65, -30, 21, 14, -83, -32, -49, -67, -22, -18, 2, 24, 42, 29, 25, 2, -78, -36, -9, 8, 0, 30, 11, -39, -35, -9, 6, 23, 22, 103, -24, 22, -75, -46, -30, -16, 4, -6, 9, 5, 51, 19, 5, -7, -33, -16, -2, -11, 27, 51, 11, 22, 1, -17, -4, 47, 44, 49, -19, -28, -12, 9, -1, -14, 9, 12, -8, 12, 27, -7, -21, -56, -39, -21, -4, 2, 17, 39, 41, -20, -18, -30, 1, 106, 61, 8, -38, -21, 23, -26, 29, 40, -18, 1, 45, 24, 16, 13, -33, -84, -53, -7, -9, -13, 19, -6, -20, -20, -6, -16, -23, 118, 62, -15, 17, -47, -16, -70, 0, -11, 0, 26, 1, 20, 13, -14, -19, -25, -12, -30, 20, 29, -6, 7, 28, 32, 20, 20, -25, 62, 10, -25, 17, -63, -96, -41, 15, 15, 12, -17, -51, -59, -20, -19, -18, -46, -40, -41, 4, 14, -2, 25, 33, 4, 13, 30, -15, 33, -10, 12, 9, -55, -60, -84, -23, 6, 72, 32, 0, -19, -109, -142, -132, -185, -207, -119, -71, -69, -81, -87, -85, -57, -51, 35, -37, 2, 17, 16, 15, 18, -26, -51, -30, -33, -20, 5, -35, -45, -91, -44, -99, -178, -192, -212, -193, -84, -76, -95, -130, -90, -78, -49, -25, -49, -10, 16, -11, -9, 16, -4, -32, -60, -59, -52, -68, -71, -100, -57, -86, -130, -98, -102, -137, -112, -103, -71, -77, -40, -52, -10, -34, -45, -7, 12, 15, 4, 2, 7, -12, -35, -31, -63, -79, -52, -29, -66, -72, -52, -18, -64, -89, -66, -40, -19, -39, -30, -21, 5, 5, 7, -10, -21, -20, 4, 20, 3, -16, 10, 2, 19, 14, 14, 4, -16, -2, -18, 4, -17, 8, 9, -20, 19, 19, -9, -8, 16, -12, 13, 9, 14, -2, 957, -16, 19, 1, -3, -1, 28, 7, 25, -4, -47, -47, -66, -39, -32, -15, -9, 3, -6, -8, -6, -10, -27, -5, -7, -13, 5, 10, 15, -19, 8, 10, -38, -7, 0, 0, -20, 43, -41, -74, -19, 13, -64, -30, -26, -32, -71, -70, -52, -52, -64, -54, -5, 0, -9, 4, -8, -20, 27, 10, 38, 17, 77, 35, 21, 32, 20, 58, 25, 53, 13, 33, 45, -6, -61, -12, -5, -27, -16, -19, 10, 5, -2, -2, -6, 20, 37, -31, -10, -47, 22, -2, -5, 16, 66, 63, 21, 35, 38, 39, 17, -12, -58, -37, -15, -28, 50, 62, 45, 25, -2, 11, 15, -10, 39, 25, -5, 3, -12, 10, 30, 30, 4, 43, 17, 43, 55, 27, 7, -25, -28, -12, -28, -26, 9, 38, -1, 7, -42, 2, 14, 16, 31, 21, -14, 41, 39, 19, 6, 20, 16, 30, 54, 66, 43, 12, -12, 11, -9, -4, -15, -32, -14, -4, 7, -36, -81, 9, 14, -8, 9, 20, -7, 24, 30, 36, 28, 34, 5, 26, 36, 27, 21, 19, 23, 4, -2, -25, -18, -13, 2, 24, 43, 17, -56, -23, -5, -9, -37, -17, -12, 7, 27, 12, 9, 31, 8, 34, 26, 12, -25, -52, 17, -10, -31, -9, -30, -62, -43, 14, 68, 40, 14, 5, -10, -32, -59, -25, 18, 11, 14, 11, 24, -1, 29, 39, 10, -82, -90, -90, -34, 1, -44, -28, -14, -44, -19, -36, 25, 56, 43, 9, -6, -14, -44, -5, 27, -11, 24, 33, 11, 27, 49, 9, -58, -135, -160, -112, -72, -18, -25, -29, -40, -31, -29, -8, -7, 3, -12, -21, -18, -19, -55, 0, -8, 34, 35, 14, -10, 26, 25, 4, -79, -122, -136, -128, -20, 23, 22, -13, 7, -9, -25, -13, -49, -23, -19, -5, -13, -20, -98, -31, 1, 26, 24, 6, 24, 0, 22, -21, -101, -111, -92, -61, -34, -20, -10, -14, 26, 16, -15, 29, 17, 3, 11, 6, 3, -24, -52, -27, 50, 44, 24, -7, -12, 0, 11, -44, -54, -91, -87, -37, -16, -9, 37, -7, -15, 26, 21, 59, 35, 6, 42, -11, 3, -22, -84, -44, 64, 48, 15, 7, 5, 7, -26, -42, -55, -67, -51, -69, -19, -8, -17, -9, 19, 19, 31, 61, 55, -23, 64, 63, 41, -23, -70, -41, 29, 31, 10, -12, -14, -20, -4, -25, -59, -74, -70, -87, -49, -18, -24, -5, 3, 24, 44, 51, 26, -33, 52, 33, 14, -26, -15, -37, 29, 47, -31, -61, -31, -3, 17, 16, -25, -72, -103, -88, -33, -9, 45, 33, 11, 23, 66, 8, -41, -58, 23, 0, 1, 27, -34, -29, -4, -54, -73, -70, -57, -25, 12, -3, -4, -77, -131, -102, -24, 35, 41, 51, 18, -12, 20, 4, -41, -62, 33, 5, 31, 24, 8, 1, -9, -121, -120, -123, -122, -130, -98, -57, -89, -141, -169, -84, 38, 73, 66, 36, 32, -24, -38, -15, -11, -25, 28, 32, 12, 37, 11, 24, 25, -76, -96, -93, -114, -146, -112, -92, -92, -121, -140, -56, 75, 105, 61, -2, 15, 0, -23, -16, -45, -38, 10, 29, 8, -27, -15, -3, 26, -26, -53, -31, -11, -30, -35, -19, -52, -85, -56, -17, 68, 74, 41, 32, 11, -2, 5, -4, -90, -70, 8, 15, 13, -15, 23, 28, 63, 31, -16, 20, 33, 71, 47, 27, 9, -26, -14, 27, 35, 61, 36, 6, 20, 47, 28, 2, -122, -75, 8, 5, -2, -20, 39, 68, 28, 51, 43, 45, 5, 45, 24, -2, -27, -38, -17, 16, 13, 9, 1, 5, 23, 24, 6, -8, -71, -83, 6, -4, 13, -8, -6, 8, 20, 31, 94, 47, -12, 10, 51, 21, -25, -20, -22, -21, 11, 10, 31, 19, 30, -2, -48, -56, -100, -65, -13, -5, -20, -4, 35, 3, 24, 33, 59, 62, 19, -5, 19, 44, 37, 15, -14, -12, 13, 16, 7, 1, -6, 6, -29, -97, -53, -17, -10, -19, -7, -14, 35, 10, 8, 9, 23, 46, 31, 66, 25, 26, 33, 37, 32, 41, 16, 4, 37, 34, -6, -45, -12, -7, 31, 37, 20, -15, -20, -20, 11, -11, -2, 45, 26, 25, 34, 64, 72, 75, 73, 81, 89, 62, 41, 21, 22, 2, 52, 69, 54, 32, 18, -7, -5, 3, -17, -8, 12, 10, -10, 26, 52, 48, 31, 41, 25, 65, 57, 44, 68, 77, 60, 33, 53, 11, 26, 36, 44, 24, 15, -8, -19, 7, -18, -7, -19, -18, 18, -14, -14, 0, -14, -6, 5, -14, 18, 4, -16, 13, 3, -8, -9, 18, 9, 5, -11, -2, -5, -19, -5, -11, -14, -1094, -9, -17, 9, -20, 18, 48, 66, 19, 58, 32, 63, 73, 110, 131, 49, 64, 36, 44, 71, 16, 27, 37, -4, -7, 8, -6, 8, -2, 17, 9, 4, 29, 39, 60, 62, 56, 14, 55, 63, 44, 56, 138, 51, 41, 59, 127, 115, 139, 142, 108, 102, 50, 7, 3, 17, -12, 9, -19, -14, -28, 1, 2, 43, 66, 31, 12, -8, -27, -7, 15, -23, 4, -9, 31, 55, 76, 30, 34, 65, 22, -17, 30, 19, -18, -15, -21, -58, -14, 69, 17, -10, 41, 6, -14, 5, -25, -1, -28, -32, -30, 5, 7, -37, -17, -16, 7, 17, 49, -25, 24, -8, -16, -7, -6, -2, 3, 63, 20, -7, 4, -15, 20, 23, 7, 0, 4, -18, -44, -11, -45, -45, -19, -21, -14, -19, -8, -46, -12, -9, 9, -8, -56, -33, -26, 4, -19, -4, -15, -14, 1, -9, 14, -13, -5, -43, -55, -46, -41, -44, -9, 9, -11, -6, -3, -20, -50, 4, -8, -4, -61, 11, 23, -32, -29, -14, -12, -4, -10, -29, 12, 6, -9, -32, -33, -50, -19, -56, -16, 17, 9, -10, -42, -36, 17, 15, -18, -7, 24, 25, 39, -6, -43, -62, -56, -10, -14, 6, 32, 1, 9, -36, -85, -80, -42, -30, 7, 11, -40, -54, -29, -65, -43, -34, -2, -18, 17, 10, -76, -56, -56, -48, -67, -9, 16, 19, 39, 4, 2, -56, -88, -72, 6, -31, -36, -23, -22, -69, -64, -60, 1, -28, 5, 3, 55, -15, -181, -166, -62, -38, -28, -6, 16, 15, -12, 25, -8, -28, -74, -4, 13, -60, -47, -38, -60, -80, -43, -39, 4, 30, 16, -56, -16, -61, -127, -159, -49, -34, -59, -2, 15, 5, 18, 2, 14, 32, 23, 11, -18, -35, -14, -49, -65, -71, -44, -25, -44, 50, 9, -3, -28, -144, -155, -93, -28, -41, -16, 10, -2, 31, -4, -2, 11, 41, 19, 17, -5, -40, 4, -3, -23, -28, 4, -41, 1, 25, 26, -4, -15, -84, -152, -80, -36, 13, -11, 25, 11, 38, -5, 12, 19, 48, 10, -11, -28, -70, -16, -48, -12, -68, 1, 20, -35, 31, -6, 11, 60, -38, -100, -56, -27, 32, 27, 51, 1, -1, 23, 41, 26, 26, -32, -61, -47, -58, -25, -19, 7, -34, 44, 39, -8, -15, -29, 45, 42, -27, -86, -41, 25, 47, 67, 49, 4, 9, 43, 25, 61, -29, -96, -94, -84, -30, -1, 19, -3, 30, 110, 36, 4, -7, 7, 46, -13, -22, -67, 46, 58, 50, 47, 45, 31, 5, -3, 30, 33, -45, -122, -112, -81, -17, 27, 37, 58, 65, 89, 62, 1, -19, 2, 67, 41, -25, -52, 17, 56, 44, 93, 21, 20, 8, -16, 6, 35, -40, -53, -29, -11, 13, 72, 65, 75, 81, 55, 25, 8, -11, -7, 66, 19, -43, -97, -2, 14, 10, 42, 5, 3, -43, -12, -5, 43, -28, -26, -12, 7, 40, 67, 71, 91, 36, 9, 16, 15, 5, -25, 8, 43, -15, -57, -43, -19, 3, 21, -8, -3, -40, -22, 40, 25, 16, 0, 8, 22, 23, 35, 77, 75, -17, -13, 2, 36, 19, -6, 34, 32, -16, -100, -52, 8, 0, -5, 30, -19, -40, 2, 20, 22, 37, -25, -8, -22, -36, 24, -21, -30, -74, -35, -4, -4, -17, -42, 6, 2, 1, -62, -50, -42, 4, -1, 27, -5, -16, 13, 61, 45, 22, 32, -9, -23, -42, -25, -45, -88, -130, -71, 21, 0, 9, 12, 16, 47, 34, -62, -58, -53, 8, 16, 5, 38, 38, 48, 50, 77, 37, 17, 11, -25, -29, -44, -63, -51, -104, -75, 59, 12, -20, -9, -12, 7, 1, -5, -36, -51, -35, -26, -4, -4, -15, -17, 2, 10, 21, 6, -28, -57, -101, -112, -26, -30, -16, -50, -14, 27, -14, -10, -9, 13, 2, -23, -15, 1, -55, -26, -27, -23, -51, -60, -49, -67, -84, -82, -92, -86, -136, -74, -77, -95, -46, 6, 46, 15, -7, 3, 17, -1, -14, 13, 27, -30, -57, -65, -58, 11, -20, -55, -43, -68, -81, -81, -128, -93, -82, -94, -94, -50, -45, -30, -12, 44, -9, -16, -20, 20, 0, -17, -36, -40, -47, -27, -92, -21, -62, -13, -2, -21, 1, -65, -76, -52, -57, -58, -33, -21, -10, -13, -20, 1, -19, 17, 16, -19, -11, 4, -64, -45, -45, -61, -22, -15, -42, -18, 35, 48, -43, -68, -52, -32, -12, -48, -47, -46, 9, -12, -11, 0, -19, 16, -13, 5, -15, -15, 2, 20, 20, 0, 19, -8, 20, -19, 10, -9, -17, -10, 6, 17, -13, -8, 6, 20, -17, -11, 16, 9, 15, -14, 2408, 15, 10, 3, 17, 6, 11, 28, 5, -6, -4, -28, -74, -70, -123, -41, -51, -34, -44, -41, -66, -38, -47, -14, 2, 4, -20, -8, 6, 10, 19, 5, 15, 32, -19, 0, -31, -48, -29, -1, -38, -24, -43, -33, -13, -45, -114, -77, -93, -124, -79, -43, -27, -8, -19, 9, 9, -14, -40, -9, 26, 47, 5, -47, -42, -28, 34, 36, 4, 59, 7, -11, -16, 16, 24, 6, -63, -50, -53, -57, -7, 12, 7, 16, 5, 9, -13, -52, -41, -24, -13, -10, 22, 12, 9, -24, 4, -6, 24, -38, -28, -2, -29, 2, -9, -7, -10, 12, -27, 11, -5, -12, 4, 16, 0, 24, -31, -40, -51, 3, 46, 16, -4, -15, 30, 19, -9, -34, -66, -65, -26, -50, -33, -79, -24, 28, 18, 29, -42, -6, 1, -25, 37, -6, -18, 2, -24, -3, 16, 15, 42, 52, 40, 9, -1, -13, -3, -13, -29, -33, -64, -77, -84, -19, 21, -33, -95, 4, 13, 15, -48, -25, -21, -40, -36, -35, -11, 9, 8, 32, 22, 16, 21, 37, 23, 34, 6, -16, -14, -65, -36, -42, 35, -37, -61, 2, -9, 27, -13, -5, -35, -55, -24, 3, 15, -12, 15, 17, 5, 9, -2, -10, 13, -2, 9, 2, 2, -60, -28, -43, 11, 15, 14, 31, 14, -15, -30, -20, -25, -61, -19, 22, 31, 10, 12, 31, 4, -11, -15, -19, 21, 48, -9, -25, 17, -22, -23, -1, 5, 47, 19, -21, 0, -41, 6, -32, -4, -13, -29, 14, 34, 50, 36, 30, 11, 23, 17, 14, 77, 50, 40, 33, 7, 26, -15, -16, -25, -17, 30, 13, -49, -45, -8, -35, 14, 51, 6, 17, 75, 49, 94, 67, 11, -4, 26, 22, 5, 15, 5, 8, 15, 39, -6, -41, -57, -24, 17, -11, -18, -51, -43, 0, 47, 18, -4, 14, 59, 69, 46, 18, -2, 10, 42, 6, 29, 21, 10, 18, 39, 63, -6, -31, -59, -3, 26, 15, -14, -35, -17, 42, 41, 75, 42, 30, 28, 33, 45, 7, 3, -38, 7, 23, 45, 22, 65, 51, 46, 7, 16, -39, -42, 17, 59, 14, 19, -13, -45, 36, 102, 108, 67, -1, -11, -6, -11, 29, -18, -19, -39, 25, 31, 66, 41, 35, 34, -4, -17, 27, -22, -7, 13, 53, 5, -18, 14, 33, 89, 100, 65, 0, -10, -12, -22, -3, 21, 21, -15, 35, 65, 42, 24, 16, -2, 32, 48, 32, 30, -14, 6, 35, 5, -65, 38, 57, 83, 75, -12, -15, -62, -44, -7, 20, 53, 3, 37, 110, 115, 50, 3, 3, 30, 31, 59, 73, 9, 41, -7, 26, 6, -32, 25, 22, 43, -19, -60, -87, -62, -36, -10, 25, 66, 29, 55, 140, 101, 40, 44, 55, 7, 24, 23, 25, 30, 21, 9, -59, 25, -64, 43, 82, 88, -39, -104, -83, -53, -56, -19, -23, -4, 16, 71, 127, 104, 62, 58, 39, 24, 34, 43, 51, 70, -16, -45, 4, -19, -32, 1, 61, 90, -11, -89, -33, -73, -55, -63, -59, -54, -39, 17, 91, 112, 93, 41, 46, 13, 39, 33, 98, 74, 10, -9, 3, -8, -15, 6, 96, 84, -15, -44, -47, -43, -89, -87, -100, -100, -53, -16, 60, 77, 64, 39, 15, 38, 47, 72, 119, 82, 32, 15, -86, -32, 29, 49, 37, 38, 38, -20, -23, -59, -44, -72, -67, -82, -71, -26, -25, 17, 41, 25, 30, 41, 75, 68, 57, 31, 49, -17, -28, -12, 16, 44, 67, 91, 83, 46, -22, 0, -31, -83, -104, -124, -92, -42, -52, -29, -5, 0, 34, 43, 43, 23, 56, 79, -8, 2, 7, -3, 29, 42, 43, 110, 105, 66, 27, 42, -18, -34, -66, -102, -79, -70, -50, -34, 25, 23, 14, 27, 8, -11, 25, 56, 34, -21, -5, 1, 11, -4, 74, 136, 135, 103, 111, 47, 20, -15, -38, -90, -101, -82, -44, -25, -2, -10, -10, -24, -13, -22, 34, 20, 18, -17, -9, 2, -6, 24, 24, 31, 45, 37, 72, 22, 10, -26, -53, -72, -47, -42, -51, -38, -35, -5, -1, 12, 25, -8, 47, 27, -32, -36, 20, 15, 4, -13, -19, -13, 3, 34, 15, 23, 27, 11, -3, -57, -27, -30, -50, -55, -23, 10, 18, 3, 40, 13, 4, -2, -36, -19, -12, 0, 11, 6, 14, -7, 7, 28, 64, 31, 25, 24, -12, -41, -34, -10, 11, 34, 22, 4, -1, 16, 12, -3, 22, 5, -16, -18, -16, 13, -3, -5, -3, 6, -2, 3, -4, 15, 20, -6, -15, 16, -15, -14, 23, 12, -8, -16, 5, -15, 8, -14, 2, -13, 19, -17, -8, -17, -560, -12, 7, -3, 14, 6, -4, -14, 14, 33, 21, 10, 36, 20, 28, 9, 9, 10, -14, -18, -6, -17, -10, -17, -4, -10, -10, -17, -15, 9, 3, -18, 7, -29, -42, -10, -7, -23, -4, 14, 6, -59, -82, -72, -29, -68, -73, -38, -71, -8, -56, -37, 42, 5, -15, 9, 16, -11, 1, -13, 29, 15, 38, 8, 5, -48, -25, -88, -115, -95, -50, -45, -32, -39, -81, -44, -73, -80, -142, -113, -82, 38, -1, 7, -13, 19, 18, -8, 5, 9, -34, -40, -60, -25, -31, -49, -50, -56, -40, -22, -26, -36, -18, 12, -18, -21, -42, 3, -55, -32, -43, -4, 1, -20, 35, 1, -23, -22, -55, -65, -53, -55, 8, 15, -4, -15, -19, 13, 21, -22, 16, 8, 8, -23, -13, 12, -34, -51, -75, 5, -11, 20, 34, 11, 22, -2, -45, -73, -25, -35, 12, 24, 6, -35, 19, 14, -24, -26, 12, 4, -12, 19, -7, 9, -32, -103, -48, -19, 24, 12, -9, -17, 2, -25, -73, -77, -61, -56, -10, 16, -19, 3, 8, -39, -34, -15, 14, -3, -4, -18, -11, -9, -52, -98, -72, -38, 21, 6, 22, -5, 13, -40, -88, -102, -47, -1, 23, 25, 29, 14, -8, -43, -49, -19, -2, 3, 4, -4, 31, -22, -77, -168, -17, 13, -3, 30, 4, -9, -10, -24, -86, -93, -71, -29, 15, -3, -10, -15, 21, 5, 10, -5, 13, 8, -7, -15, -19, -31, -18, -124, -19, -35, -4, 20, 33, 8, -21, -44, -48, -54, -66, 0, 15, -3, -16, 4, 30, 4, -15, 12, 16, 4, 8, -7, -27, -20, 43, -18, -43, 6, -29, -57, -49, -43, -12, 20, -5, -32, 27, 14, 13, -18, -39, -12, 20, 3, -21, -5, 30, 7, 8, 1, 2, 47, 43, -1, -81, 17, 18, -47, -47, -81, -21, -9, -33, -42, 3, -25, 11, -37, -42, 2, 40, 9, 1, -5, -18, -45, -47, -48, -6, 68, 19, -2, -33, -8, -14, -44, -90, -57, -83, -31, -55, -63, -16, -29, -13, -37, -3, 6, 17, 3, 32, -25, -37, -33, -16, -9, -18, -1, -16, 9, 9, 4, 21, -33, -56, -56, -89, -142, -116, -111, -28, -56, -68, -43, 27, 20, 14, 31, 2, -34, -23, 5, -15, -58, -89, -78, -37, 40, -9, 6, 8, -6, -77, -105, -133, -129, -156, -136, -82, -75, -74, -3, 18, 23, 34, 41, 26, 0, -22, -17, -43, -68, -122, -92, 2, 8, -40, -14, 13, -24, -8, -49, -43, -74, -69, -57, -65, -50, -36, 28, 16, 48, 35, 41, 67, 4, -89, -110, -128, -96, -80, -11, 50, -27, 4, 4, 15, -34, -11, 60, 73, 58, -3, 17, -69, -44, -11, 31, 34, 50, 29, 106, 71, -49, -164, -188, -187, -172, -90, -8, 49, -45, 6, 21, 4, -42, -7, 56, 68, 30, 26, -13, -55, -5, -6, 27, 55, 78, 110, 126, 86, -67, -164, -207, -152, -120, -97, -40, 10, -18, -31, -2, -49, -24, 2, -37, -20, -43, -19, -30, -59, -10, 7, -20, 29, 45, 116, 117, 31, -56, -155, -180, -193, -121, -79, -10, 30, -67, -44, -20, -41, 8, -28, -19, -27, -9, -34, -31, -59, -36, -13, -11, -39, 2, 83, 84, 12, -41, -166, -161, -117, -110, -95, -10, 22, -35, -31, -79, -6, 7, 46, -51, -42, 49, 17, 16, -8, 4, -26, -18, -2, 12, 21, 33, 22, -47, -110, -173, -128, -91, -110, -43, 32, -28, -27, -66, -1, 26, 56, 10, 13, 74, 13, 24, 45, -19, -30, -13, -44, -25, -9, -41, -57, -64, -110, -156, -135, -121, -59, -34, 11, 12, -68, -34, -20, 5, -4, -51, 2, 52, 22, 38, 0, -15, -41, 1, -33, -22, -47, -91, -127, -124, -135, -123, -150, -79, -22, 20, 6, 11, 19, 18, 18, -42, -18, -54, 1, 116, -6, 36, -28, -2, -19, -5, -32, -49, -59, -88, -150, -123, -94, -78, -70, -78, -29, -23, 38, 9, 4, 1, 5, -7, -1, -21, -17, 5, 16, 2, -30, -67, -34, -37, -74, -51, -104, -149, -146, -164, -122, -98, -95, -10, -41, 14, 52, 19, 6, -5, -4, -12, -19, -19, -8, -4, 71, 54, 59, 101, -14, -30, 0, -23, -12, -62, -106, -67, -63, -62, -52, -22, 6, -22, 23, -9, -18, -8, 10, -1, -2, -18, 10, -14, 36, 29, 52, 34, 40, -49, -34, 3, 19, -27, -38, -52, -1, -20, -3, -20, -6, 18, -17, 7, -1, -16, 6, 2, 8, 0, 7, -8, 20, -15, 16, 10, -1, -18, 4, 19, 2, -8, 18, 3, -14, 17, -20, 8, 14, -12, 3, 6, 7, -11, -3, 814, -19, 16, 1, -12, 45, 34, -1, -4, -5, 3, 26, 21, -21, -22, 51, 16, 10, 39, 39, 18, 17, 16, 61, 24, 1, 14, -19, -3, -1, 10, 17, -22, -4, 91, 47, 33, 87, 34, 13, 56, 54, -37, 27, -15, 4, -17, -22, 0, -5, -39, -38, -69, 1, 2, 15, 12, -18, -16, 10, 36, 31, 86, 39, 33, 106, 74, 39, 61, 33, 31, 30, 64, 52, 31, 54, 60, 52, 20, 53, 50, 22, 0, -13, 4, -13, 15, -45, 24, -29, 21, 51, 4, 50, 37, 55, 23, 28, 37, 24, 23, 16, 54, 48, 22, 23, 54, 71, 76, 58, 17, 19, -10, 10, 13, -43, -4, -34, 8, 9, 23, 15, 15, 53, 17, 36, -3, -32, -3, 32, 59, 24, -23, 17, 33, 38, 53, 63, 34, -15, 0, -6, -7, -73, -51, 31, 25, 1, -12, 24, 55, 40, 7, 34, -9, -24, 5, -12, -27, -2, 8, -6, 0, -16, -25, 12, 8, 9, 6, 20, 4, -66, 2, 53, 40, 2, -14, 27, 11, 22, -23, -28, 7, -3, -11, 10, -17, -23, -17, 1, -6, -5, 3, -13, -22, 0, -20, 29, -18, -64, 3, 50, 22, -29, -40, -22, 11, -1, -29, -18, -17, -19, -1, -9, -32, -21, -26, -17, -1, -7, -19, 18, 34, 32, 17, 9, -12, -10, 24, 10, -2, -2, -24, -34, 14, 26, -9, -9, -16, -25, -28, -92, -78, -87, -65, -29, -31, -21, 5, 34, 69, 47, -12, -14, -12, -34, 0, 3, 28, 21, 14, -41, 10, -3, -19, -10, -44, -78, -74, -67, -131, -126, -79, -67, -28, -12, -20, 34, 24, 4, 36, 34, -5, -46, 26, 50, 2, -8, -19, 0, -7, -2, -35, -54, -44, -66, -88, -97, -77, -104, -82, -83, -47, -18, 4, 20, -1, 23, -4, 12, 6, -38, 100, 54, 26, 1, -27, -6, -44, -47, -67, -32, -85, -93, -78, -62, -37, -29, -21, -22, -41, -9, -24, 13, 14, 27, 7, -22, 25, -15, 108, 63, -15, -25, -29, -57, -25, -50, -46, -57, -101, -113, -82, -54, 11, 14, 22, 33, 13, 8, -18, 24, 52, 0, 37, 2, -32, -62, 101, 76, -38, -48, -68, -64, -59, -53, -58, -60, -90, -116, -51, -3, 36, 33, 33, 12, 29, 28, -32, 12, 73, 16, 13, -50, 22, 6, 39, -46, -62, -71, -55, -74, -15, -24, -69, -101, -55, -63, 20, 59, 83, 66, 41, 42, 49, 22, -30, -1, 76, 2, -4, -41, 55, 56, -9, -47, -76, -63, -65, -50, -5, 11, -18, -53, -44, 16, 67, 101, 99, 74, 36, 45, -5, 5, -6, 20, 49, 28, 21, -10, 86, 101, 39, 9, -23, -25, -12, 36, 46, 27, -34, -9, -2, 74, 84, 94, 59, 34, 16, -34, -25, 2, 29, 83, 74, 37, 31, 11, 69, 123, 95, 65, 18, 39, 56, 37, 50, 27, 7, 21, 46, 125, 78, 70, 71, 47, 8, -15, 10, 5, 22, 64, 70, 36, 45, 43, 18, 129, 93, 48, 50, 14, 4, 32, 56, 19, 7, 25, 37, 55, 60, 31, -10, 6, -19, -13, 15, 19, 30, 5, 4, 62, 38, -6, -24, 67, 93, 77, 55, 35, 8, -24, -14, -22, -3, -4, -9, 14, 39, 17, -17, -2, -4, 22, -12, 0, -29, -9, 0, 45, 26, 56, 15, 22, 11, 21, 15, 14, 13, -17, -28, -19, -33, -50, -46, -16, -22, -2, -30, -18, -17, 37, 8, -6, 20, 52, 31, 68, -16, 27, 55, 73, 37, -18, -8, -15, -33, -26, -35, -37, -69, -44, -29, -16, -20, -21, -53, -65, -40, -1, 10, 44, 71, 45, 18, 20, 5, 1, 41, 48, 24, 18, -32, -33, -59, -52, -51, -58, -52, -63, -11, -29, -30, -36, -45, -4, 27, 45, 31, 61, -3, 32, -10, 6, -10, -58, 33, 17, -9, -41, -28, -38, -69, -32, -16, 4, -18, -6, -42, -32, 2, 10, -4, 0, -36, -6, -28, -15, -14, 41, 2, 12, 11, -19, 45, 5, -22, -41, -19, 5, -8, -11, -2, -13, -14, -22, -48, -34, 14, -24, -46, -20, 6, -26, 14, 6, -22, 14, -14, -6, -11, -5, 9, -1, -1, 15, -29, -19, -12, -14, -3, -32, -29, -60, -98, -106, -63, -55, -30, -18, -31, -3, -43, -9, 14, 23, -3, 16, -19, 9, 5, -10, 2, 24, -1, 0, -13, -3, -27, 11, -3, -37, -11, 8, 10, 23, 12, -21, 26, 35, 11, -3, 14, 10, -19, -18, -1, 11, -2, -17, 14, 7, 17, -9, 3, 13, -15, -5, 0, 0, -20, 1, -19, 19, 4, -13, 5, -4, 3, 4, -8, -18, -19, 13, -12, 40, 16, 5, 18, 6, 15, -18, -24, -35, -19, -12, -60, -72, -45, -148, -104, -88, -65, -85, -81, -40, -29, -34, 7, 24, -20, -20, 17, 15, -1, -12, 0, 7, -19, -49, -62, -69, -99, -101, -150, -86, -56, -115, -127, -105, -108, -95, -100, -127, -70, 46, 64, 17, -7, -18, -1, -3, 2, -6, 4, 18, 73, 59, 33, -11, -72, -46, -68, -84, -76, -41, -45, -51, -27, -17, -18, -18, -16, 4, 68, 77, 71, 1, 20, -15, -20, 7, -9, -19, 40, 49, 0, 6, 3, -10, -4, -34, -50, -10, -19, -37, -8, 62, 82, 43, 66, 116, 148, 127, 90, 15, -12, 6, 16, 62, 23, 19, 2, -18, -14, -27, 4, 2, -24, -41, -50, -17, -38, 25, 39, 107, 81, 89, 100, 105, 150, 106, 55, 37, -3, -5, 8, 55, -21, 8, -25, -26, -24, -47, 12, -18, -24, -38, -60, -60, -50, -16, 56, 66, 55, 84, 57, 87, 85, 120, 77, 42, -16, -16, -4, 4, 2, -24, -45, -31, -16, -43, -31, -33, -34, -59, -91, -75, -45, -35, 25, 49, 68, 72, 57, 19, 57, 64, 93, 51, 9, 11, -5, 1, -35, -55, -68, -63, -65, -78, -43, -36, -56, -56, -77, -51, -34, -33, -6, -32, -23, -6, -34, -5, 14, 3, 65, -2, 18, 15, 10, -24, -13, -81, -148, -152, -56, -67, -71, -57, -70, -33, -26, -19, -53, -63, -71, -111, -166, -156, -119, -97, -55, -22, 48, 5, -27, 22, -26, 47, 2, -31, -92, -119, -55, -82, -44, -40, -43, -23, -10, -46, -59, -56, -60, -158, -200, -249, -208, -150, -127, -47, -19, -28, 14, -29, -54, -5, -22, -70, -62, -113, -53, -49, -43, 10, -15, 11, -23, -31, -55, -74, -101, -79, -130, -185, -201, -168, -141, -58, -22, -37, 21, 0, -56, -66, -90, -85, -106, -76, -32, -6, -11, 24, 6, -14, 37, 5, 16, 9, -16, -28, -54, -48, -86, -129, -76, -47, -35, -40, 18, 0, -30, -31, -89, -111, -31, -61, 22, 8, 2, 39, 25, 34, 72, 44, 29, 55, 32, 45, 54, 9, -40, -62, -47, -34, -5, 36, 56, 3, -34, -79, -95, -71, -39, -30, -13, 19, 42, 16, 50, 52, 57, 40, 53, 51, 47, 33, 55, 55, 42, -29, 30, -52, -42, 0, 37, 5, -47, -86, -39, -35, -31, -6, 35, 50, 57, 11, 27, 56, 83, 46, 50, 48, 10, 54, 27, 39, 33, -2, -24, -60, -94, -46, 18, 17, -24, -19, -15, -16, -30, -30, 24, -5, 15, 14, -17, 56, 56, 58, 44, 33, 35, 39, 16, 24, 11, -10, -98, -124, -76, -8, 1, -18, -54, 21, 33, -27, -34, -12, 9, 1, 2, 1, -14, 31, 35, -20, -44, -10, -15, -5, 10, 46, 8, -34, -76, -52, -46, -34, -15, -9, 2, 39, 63, 0, -33, -18, -6, 34, 12, -24, 12, 23, 37, -51, -67, -34, -46, -34, 14, 29, -3, -73, -56, -14, -3, -6, -30, -4, 13, -2, 13, 48, -16, 8, 20, -2, 2, 12, 27, 37, -18, -39, -27, -14, -4, -2, 54, 44, -5, -28, -33, -25, -31, -9, -7, -29, -15, -16, 73, 66, 14, 1, 31, 19, -7, 6, -9, -18, -41, -70, -69, -35, 7, 34, 45, 7, -16, -1, -20, -16, -15, 19, -34, -11, 18, 12, 4, 18, 16, -13, -18, -7, -18, -34, 8, -39, -54, -39, -19, 11, 20, 16, 24, 7, -19, -36, 26, -20, -39, 20, -53, 2, -5, 23, -32, 25, 9, 33, -15, -26, -30, -30, -27, -55, -67, 0, 7, -19, 25, 34, 33, 1, -21, -38, 10, -21, -25, 28, -13, -12, -14, -31, -37, 16, 41, -33, -49, -55, -77, -80, -21, -11, -23, -46, -23, 1, 2, 39, 58, 23, -39, -19, 4, -19, -47, -28, 14, 0, -21, -27, -46, 6, 25, 23, 18, -4, -6, -67, -83, -69, -63, -103, -38, -4, -38, -44, -85, -75, -18, -27, 36, 22, 26, 1, -10, 18, 11, 10, -58, -61, -36, -5, 0, -3, 0, -39, -86, -109, -93, -58, -95, -20, -5, -68, -81, -34, -48, -10, 3, 33, 17, -10, -14, 12, -20, 1, 1, 0, -34, -34, -26, -4, 51, -26, -11, -54, -38, -57, -53, -29, -29, -82, -42, -13, -27, -30, -4, -26, 3, 8, 14, -10, 13, -9, -1, -7, -18, -42, -34, -20, -5, -8, -45, -55, -36, -29, -41, -25, -16, -9, 4, -30, -23, -14, 13, -20, 12, 6, -8, -9, 15, -1, 1, 20, 16, 3, -8, -8, 4, 12, 5, 7, 8, -22, -27, -5, -19, -12, -7, -14, -12, 7, 19, 18, -19, -20, -10, -14, -772, -2, 4, 4, -2, 5, 5, 21, -18, 11, 37, 47, 38, 27, 63, 17, 28, 18, 74, 15, 46, 38, 28, 22, 4, 1, 4, 13, 12, -12, -2, -2, 17, -2, 59, 65, 36, 68, 47, 55, 86, 73, 86, 69, 35, 8, 47, 38, 7, 4, 44, 15, 26, -6, 16, 11, -1, 17, -2, 7, 38, 53, 37, 19, -18, -21, -34, -16, 9, -2, 12, 28, 54, 42, 15, 43, 63, 34, 67, 113, 46, 35, -7, -20, 6, 4, 45, -40, -72, -44, -53, -37, -55, -91, -55, -2, -31, 10, 12, 1, -7, 25, 37, 42, 1, 13, 59, 76, 91, 90, -1, 4, 5, -9, 42, -70, -33, -53, -69, -80, -36, -27, -6, 19, -1, 52, 14, 19, 28, 32, 61, -9, 1, -3, 48, 77, 118, 72, 21, 5, 5, -15, 9, -57, -65, -41, -13, -41, 16, 15, 6, -1, -3, 35, 20, 27, 49, 68, 67, 53, 45, -7, 15, 57, 51, 42, -39, -3, 11, 7, -18, -16, -43, -27, -20, -3, 0, 32, 27, -4, 25, 7, 21, 36, 45, 42, 72, 60, 81, 84, 29, 55, 60, 35, -11, 4, -4, 15, -9, -17, -4, -22, -8, -17, 5, 13, 0, 21, -4, 25, 11, -31, -49, -30, 5, 27, 39, 13, 22, 35, 27, 38, 9, 20, 13, -5, -54, 13, -31, 1, -15, 10, 21, 8, -2, 5, 4, 13, 2, -98, -139, -161, -118, -72, -53, -36, -11, -27, -14, 57, 50, 19, -12, -1, 15, -31, -97, -67, -1, 33, -13, -20, -18, -8, -1, 6, -36, -165, -245, -236, -275, -263, -157, -109, -102, -101, -45, 47, 37, 31, 41, -7, 16, -85, -15, -20, -43, -10, -15, -5, -11, -5, -35, -20, -57, -81, -103, -143, -218, -246, -250, -206, -140, -94, -84, 10, 13, 40, -3, -17, -117, -128, -9, 9, 13, 11, -7, -16, 23, -17, -42, -12, -2, 0, 24, 32, -34, -99, -151, -156, -127, -66, -36, -17, 29, 49, 11, -19, 2, -94, 3, 52, 58, 43, 22, -10, -14, -11, -37, -9, -6, 35, 33, 18, 41, 8, -79, -118, -93, -80, -43, -4, 12, 20, -4, -41, -79, -61, -12, 18, 23, 47, -16, -55, -36, -45, -5, 3, 8, 24, 8, 2, 25, 4, -31, -59, -27, -61, 13, -22, 28, -8, 22, -19, -19, -53, -58, -63, -13, -17, -6, -60, -51, -14, -24, -19, 30, 20, 25, -18, -2, -7, 10, 6, 4, 30, 49, -9, 10, -2, -17, 44, 77, -41, -135, -61, -8, -8, -15, -48, -30, -7, -22, -15, 24, -22, 6, -1, 14, 0, -3, 26, 13, 28, 65, 16, -1, -9, 2, 21, 59, 65, -2, -30, -4, -1, -16, -18, 15, 19, -22, -32, -20, 19, 20, 3, -14, -47, 11, 31, -5, 2, 62, 41, 41, -29, 1, 37, 81, 102, 17, -63, 7, 19, -19, -35, -26, -26, -42, -34, 9, 22, 38, -6, 3, -2, 35, 31, 15, 18, 39, 90, 5, -4, 22, 57, 0, 41, 24, -40, -9, -3, -37, -55, -23, -42, -34, 40, 40, 33, 25, -7, -5, 1, 42, 31, 19, -12, 33, 2, -1, 2, 10, 12, -7, 20, -5, -39, -25, -14, -10, -7, 2, -11, -22, 32, 49, 36, 30, 31, -12, -3, 4, -26, -1, 4, -18, 25, -13, 10, 10, 53, 5, 10, 3, -46, -6, 23, 18, -7, -9, 10, 4, -17, 26, 44, 41, 32, 19, 11, 13, -18, -7, -15, 26, 21, -12, -13, -4, 20, 23, 53, 16, 8, -22, -29, 4, 0, 0, -5, -2, 3, 31, 14, 14, 17, 29, 8, 10, -10, -4, 17, 54, 30, 19, -11, 16, -18, 5, 53, 16, 44, 32, -42, 6, -31, -27, -17, 4, 18, 11, 18, -22, -22, -23, -11, -12, -16, 40, 64, 10, 20, 30, 15, 18, -54, -11, 33, 19, 21, 55, 16, -39, -19, -17, -52, -40, 15, -8, 10, 5, 21, -14, -21, -22, 6, 9, 61, 56, 36, 21, 24, -10, 6, -16, -50, 18, -28, -16, -18, 14, -5, -14, 13, 28, 71, 16, 8, 22, -33, -15, -3, -11, -7, -21, -20, -17, -3, 9, -20, 16, 0, -14, -4, -29, 9, 4, 2, 18, 37, 34, 49, 63, 67, 24, -34, -43, -67, -36, -61, -47, -23, -21, 10, -21, -4, -20, 18, 16, -11, -19, -20, 13, -15, 6, 0, -20, 14, -4, -25, -5, 13, 34, -24, -32, -26, -1, 0, -36, -17, -1, 2, 1, 21, 18, -1, 2, 6, 10, -17, 10, 18, -13, 11, -11, -3, -16, 5, 2, 21, 14, -5, -5, -13, -5, -2, -9, -8, -20, -14, -1, -4, 1, -17, -7, -114, -3, -3, 13, 18, 34, 41, 41, 17, 20, 23, 73, 59, 48, 69, 23, -11, -2, 28, -8, 28, 27, -10, -15, 3, 16, -8, 5, -5, 8, -6, -4, 13, 35, 31, 55, 23, -34, 32, 97, 60, 42, 45, 64, 80, 82, 105, 108, 96, 39, 36, 32, 7, -3, -17, -18, 4, -3, -34, -17, -15, 20, 9, 19, -3, 12, 3, -45, 19, 1, 9, 70, 85, 111, 179, 159, 76, 79, 112, 108, 68, 23, 36, 12, -11, -17, -35, -74, -97, -42, -85, -27, -22, -64, -120, -69, -14, -36, -5, 2, -51, -12, 7, -17, 16, 30, 31, 32, 51, 61, 64, -6, 0, 20, -20, -13, -43, -79, -68, -52, -23, -55, -19, -46, -14, -6, -38, -41, -60, -45, -35, -52, -37, 7, -49, -32, -13, -16, 20, 14, 20, 6, 16, -33, -40, -63, -46, -35, -30, -25, -54, -23, -40, -40, -62, -45, -33, -48, -54, -79, -55, -9, -29, -67, -67, -39, -38, 20, -7, -15, -54, -70, -97, -52, -34, -25, -49, -55, -47, -48, -63, -61, -86, -37, -58, -79, -74, -51, -11, -19, -17, -56, -36, -30, -5, -10, 1, -4, -36, -85, -29, -30, -36, -37, -36, -27, -65, -87, -89, -44, -23, -57, -83, -61, -32, -16, -29, -14, -4, -14, -39, -11, -29, 15, 14, -61, -55, -89, -9, 9, -26, -12, -30, -34, 5, -33, 11, 7, -4, -27, -12, -28, 21, -15, 2, -12, -18, 29, 14, 31, -11, -14, 12, -45, 6, -69, -26, -32, -9, -8, -26, 29, 48, 70, 59, 72, 23, 2, 32, 62, 16, 18, 17, -3, 20, 37, 47, 42, 54, -1, 23, -55, -25, -56, 24, 7, -8, -21, 7, 75, 100, 99, 57, 30, 16, -13, 33, 54, -11, 21, 51, 30, 33, 2, 9, 24, 45, 48, 17, -72, -101, -16, 47, 12, 45, -3, 36, 114, 123, 89, 67, 44, -11, 25, 49, 71, 54, 34, 30, 17, 31, -8, 12, 6, 42, 22, -18, -49, -57, 14, 36, 84, 90, -13, 50, 98, 86, 103, 38, 59, 35, 18, 68, 125, 82, 5, -9, 5, 72, -2, 8, 5, 28, 19, -5, -47, -48, 29, 54, 75, 54, 24, 43, 103, 80, 76, 58, 44, 42, 78, 91, 149, 91, 32, 13, 15, 63, 21, 4, -6, 30, 38, -11, -13, 5, 38, 55, 54, 15, 33, 64, 79, 56, 57, 69, 76, 49, 109, 122, 137, 50, 4, 3, 7, 36, 40, 4, 0, 8, -2, 0, 13, 4, 33, 21, 72, 55, 39, 57, 59, 67, 40, 80, 96, 77, 141, 94, 98, 59, -13, -21, 20, 18, 15, -1, 47, 47, 14, 31, 22, 13, 5, -21, 24, 37, 14, 41, 40, 50, 67, 51, 71, 59, 91, 85, 53, 35, 27, -25, 5, -21, 3, 12, 78, 36, -1, 33, 2, -38, -5, -14, 21, 31, 9, 39, 14, 18, 10, 9, 9, 21, 16, 0, 14, -1, -14, -6, 13, -7, -10, -4, 29, 20, 18, 17, 0, 5, -32, -52, -1, 13, 25, 6, -26, -10, 0, -19, -5, 7, 2, 2, -6, -15, 2, -28, 7, 5, -4, 6, 52, 17, 44, -5, 44, 2, -5, -52, -53, 0, -28, -9, 4, -17, -18, -5, -49, -61, -46, -21, -3, -3, -24, 6, -13, -6, -9, -10, 27, 6, 33, -26, 10, 27, -20, -18, -34, -34, -32, -12, -28, -26, -25, -26, -30, -43, -39, -54, -39, -33, -24, -28, -26, -22, -4, 24, 47, 27, 32, -3, 1, -8, 34, -41, -23, -37, -57, -26, -23, -11, 9, -6, -3, -50, -28, -41, -19, -1, -3, -9, -9, -13, 49, 39, 54, 49, 0, -11, 17, 33, 38, -35, -45, -53, -69, 5, -4, -20, 20, 9, 24, 7, 6, 14, -14, 25, 24, -9, 35, 51, 103, 60, 16, -51, 4, -4, 7, 45, 64, 37, 19, 16, -3, -2, 10, -4, -34, -2, 3, 13, 17, 12, 44, 38, 18, 37, 5, 23, 39, 45, 30, -10, -2, 13, 12, 13, 32, -4, 58, 52, 58, 89, 14, 25, -5, -60, -33, -19, -1, 33, 28, 5, 16, 24, 24, 46, 25, 34, 15, -1, 19, -2, 5, -5, -20, -20, -8, 29, 3, 39, 75, 23, -23, -33, -21, -54, -48, -5, 20, 9, -44, -49, -18, -26, -17, -8, 2, 7, 19, 7, 13, 7, -20, 17, -1, -39, -14, -3, -2, -7, -25, -35, 6, 4, -19, -18, -38, -4, -18, -12, -14, -14, 12, 0, -11, 6, -13, 17, 18, 4, -3, -9, -1, 18, 7, -14, -7, 13, -20, -13, -2, -26, -25, -1, -16, 12, -13, -3, 19, 7, -12, -17, -5, 16, -3, -17, 85, 20, 5, -3, 16, -21, -68, -46, -64, -45, -81, -126, -110, -104, -129, -50, -23, -15, -37, -59, -35, -25, -40, -2, -5, 10, -6, 0, 13, 9, -15, -8, -16, -32, -45, -75, -78, -61, -58, -38, -25, -71, -135, -90, -50, -36, -93, -147, -120, -106, -105, -81, -39, -25, -2, 9, 20, -18, 16, 2, 15, 1, -27, -41, -41, -26, -24, -38, -12, -11, -39, -9, 18, -38, -47, -48, -58, -97, -87, -104, -78, -37, 6, -4, 9, -12, -10, 22, 2, -23, -56, -66, -65, -22, -10, 10, 9, -12, 37, 36, 10, -4, -22, 42, -5, -66, -81, -54, -57, 49, -6, 4, -4, -19, 36, 26, -27, -4, -24, -34, -24, 12, 26, 39, 3, 10, -4, 29, 5, 19, 50, 70, 54, -30, -2, -9, 37, 89, 56, 19, 12, 6, 52, 20, -7, 18, 37, -9, 4, 22, 63, 41, 11, 24, 2, 31, 30, 62, 24, 41, 22, 38, 8, 27, 28, 90, 27, -17, -7, -7, 43, -2, -17, 38, 76, 24, 40, 40, 54, 63, 29, 28, 1, -3, 46, 60, 30, 45, 32, 92, 83, 32, 73, 115, 54, 23, 1, -6, 13, -29, 2, 55, 90, 81, 62, 41, 52, 52, 25, 26, -18, 20, 32, 44, 42, 82, 85, 135, 123, 65, 59, 116, 63, 42, -3, -23, 13, 24, 101, 138, 130, 41, 57, 25, 63, 68, 36, -6, -34, -12, 16, 32, 37, 53, 52, 72, 75, 55, 5, 51, -3, 15, 8, -20, -22, 25, 167, 171, 69, 39, 39, 14, 18, 29, 44, 0, -23, -32, -32, 9, 48, 40, 66, 35, 61, 33, 36, 44, 30, 6, -59, 36, 57, 51, 118, 108, 51, 10, 45, 22, -19, 18, -16, -16, -43, -49, 0, 7, 20, 23, -18, 21, 5, 31, 13, 45, 54, 16, 20, 32, 77, 190, 121, 62, -20, -13, -2, 15, -2, -32, -23, 0, 12, -10, 24, 51, 28, 40, -8, -1, -36, 6, -18, 21, 45, 14, -4, 9, 76, 138, 175, 10, -18, -41, -29, -40, -48, -52, 4, -33, 22, 25, 26, 20, 39, 22, 6, 10, -13, -10, -34, -32, 36, 3, 19, 12, 60, 61, 124, 4, -41, -58, -47, -30, -43, -15, -26, -9, 5, 21, 81, 73, 18, -4, -23, -5, -35, -24, -52, -6, -38, -29, 21, 21, 10, 23, 69, 51, -10, -36, -50, -4, 17, -20, -12, -48, -24, 42, 81, 46, -11, -17, -43, -54, -46, -39, -32, 27, -54, -8, 1, -28, 13, 34, 115, -6, -28, -50, -19, -27, -20, -18, -42, -51, -4, 67, 77, 37, -18, -36, -84, -71, -66, -23, -26, 58, -30, -46, -19, -50, 31, 50, 94, 23, -55, -73, -46, 2, 12, 11, -21, -16, -31, -4, 1, -17, -42, -74, -65, -72, -72, -12, 39, 26, -40, 12, -12, -46, 48, 24, 64, 19, -38, -28, -38, -5, -1, 23, -14, -14, -40, 1, -10, -24, -15, -36, -19, -32, -25, 22, 55, 16, -6, -77, -11, -22, -35, 27, 35, 22, -22, -17, -2, 36, 27, 30, 32, -37, -40, -35, -46, -15, 1, -15, -32, 0, -32, -1, 19, 15, 14, -61, -1, 16, -23, -7, -12, 8, -13, -15, 11, 29, 16, -4, 17, -38, -24, -30, 2, -10, 11, 21, -41, 31, -17, 28, 29, 9, -20, -58, 40, 11, -32, 5, 31, -19, -24, 4, -54, -31, -33, -28, -38, -38, -38, -42, -44, 10, -3, 18, 14, 12, 4, 50, 3, -52, -70, -15, -18, 13, -27, 37, 46, 33, 19, 2, 1, -22, -27, -59, -61, -41, -30, -33, -20, -15, -24, 10, 7, -7, -1, 12, 23, -35, 6, 32, -18, 23, 41, -16, 11, 54, 138, 90, 60, 28, 0, 30, 38, 39, 31, 20, 17, 4, 29, 46, -26, 12, 3, -9, 49, -2, 27, 1, -14, 27, 31, 35, 5, 24, 36, 49, 131, 127, 119, 165, 156, 177, 172, 171, 167, 161, 181, 180, 121, 95, 97, 33, 31, -11, -19, 15, -2, -11, 17, 37, 5, -8, -4, 35, 83, 47, 36, 70, 178, 198, 182, 208, 166, 144, 103, 116, 120, 116, 54, 36, 42, 13, -22, -8, -8, 4, -3, 7, 26, 46, 49, 27, 78, 111, 62, 53, 125, 123, 120, 109, 112, 97, 65, 83, 100, 92, 30, 21, 47, 43, -14, -10, -14, -12, 1, -13, -1, 36, 36, 43, 79, 40, 67, 53, 75, 33, 8, 74, 78, 55, 67, 25, 42, 50, 47, 15, 15, -17, 16, 7, -7, 20, -2, -18, 13, -8, 19, 11, 0, -1, -2, -14, 18, 12, 12, -6, 24, -19, 2, -3, -20, 17, 20, 5, 4, 12, 7, -6, 7, -1094, -1, -20, -15, 19, 34, -11, -26, -21, -19, 4, 45, 69, 105, 12, 87, 96, 85, 76, 40, 51, 57, 25, 34, 24, 9, -12, -3, 5, 16, 21, 14, -17, -57, -22, -44, -71, -29, -17, -26, 1, 90, 101, 64, 19, 38, 46, 21, 62, 21, -54, -67, -36, 7, 13, 10, -8, -8, 21, 20, -39, -56, -110, -48, -39, -102, -100, -18, 57, 64, -3, -24, 37, 31, 35, 44, 76, 60, 45, 12, 16, 9, -37, -13, -1, -1, 13, 53, 97, 5, 7, 16, -26, -35, -31, -16, -55, 6, -2, 0, -4, 8, -25, 1, 18, 24, -18, -6, -1, -76, 7, 4, -7, -6, -3, 0, 5, 22, 46, 71, 37, 34, 18, -5, -1, 7, 11, 25, 15, 4, 3, 12, 9, 12, 25, -5, -1, -61, -10, 8, 12, 8, -3, 11, 19, 21, 62, 59, 21, 35, 32, 23, 4, 17, 38, 14, 24, 7, 5, -11, 9, -20, -6, 49, 13, 22, 48, -5, -25, 8, 8, 23, -23, 47, -1, -15, -13, 49, 9, 7, 20, 21, 54, 43, 51, -5, -20, -5, -12, -27, -34, 29, 15, -8, 21, -2, 5, -18, 11, 30, -23, 1, -38, -29, -26, -15, -4, -28, -8, 10, 29, 66, 35, 44, 4, -29, 5, -18, 4, 17, 27, 15, 3, -51, -7, 44, 55, 59, -29, -29, -30, -28, -35, -38, -36, -29, -11, -16, 31, 47, 72, 59, 21, 30, 35, 37, 28, 35, 35, 35, -23, -22, -7, 45, 19, 50, 26, 14, 12, -39, -76, 2, -16, -3, -37, -37, -16, 22, 73, 45, 33, 4, 30, 83, -6, 1, 13, 50, -60, -9, 0, 64, 44, 80, 13, 2, -37, -73, -52, -36, -43, -37, -47, -26, -26, 9, 41, 68, 50, 81, 33, 28, 14, -26, -46, 4, -46, -30, 8, 50, 71, 64, 47, 21, -29, -11, -28, -9, -27, -29, -22, -51, -4, 5, 37, 86, 79, 67, 14, -42, -57, -86, -137, -69, -61, -38, 17, 40, 82, 77, 66, 2, 14, 37, 3, -7, -9, -19, -22, -31, -7, 31, 48, 84, 65, -31, -65, -100, -159, -192, -183, -83, -62, -7, -11, 60, 128, 97, 42, 3, 18, -1, -30, -14, -8, -44, -33, -52, -36, 38, 36, 38, -62, -160, -235, -209, -200, -215, -154, -89, 18, -29, -14, 31, 76, 84, 48, 10, 12, -16, -24, -23, -30, -37, -10, -20, -27, 21, -27, -149, -211, -254, -232, -258, -181, -123, -128, -68, 57, 32, 12, 26, -19, 37, 0, -62, -42, -7, -33, -26, -9, -36, -25, -30, -83, -120, -154, -216, -249, -181, -110, -84, -43, 23, -22, -65, -23, 7, -13, -42, -67, -34, -30, -45, -15, -23, -46, -36, -19, -16, -20, -66, -139, -175, -156, -114, -69, -46, 22, 15, 45, 69, -34, -72, -13, 14, 6, -9, -22, -11, -21, -29, -25, -32, -45, -39, -13, 4, -55, -94, -114, -106, -62, -39, 7, 50, 34, 47, 62, 56, -62, -45, 28, -27, 11, 22, -12, -59, -85, 35, 6, -42, -35, -9, 5, 14, -54, -28, -30, -4, 6, 31, 32, 47, 35, 23, 25, 47, 7, -33, -3, -3, 28, -17, -59, -121, -94, 12, 35, 20, -2, -8, -35, 22, 18, 2, 55, 34, 21, 47, 48, 17, 33, -4, 1, -2, -11, -21, 2, 33, -3, 18, -3, -94, -32, -37, 27, 16, 25, -5, -19, -6, 31, 16, 44, 59, 11, 29, 26, 32, 20, 28, 14, 15, -10, 1, 12, 15, 14, 18, -3, -93, -46, -43, -17, -1, 4, -22, -11, -6, 28, 35, 32, 15, 31, 6, 41, -7, -6, 13, 32, -13, -7, -35, 8, -5, 6, 15, 14, -3, -14, -30, -34, -30, -18, -39, -10, -10, 26, -24, -10, 21, 9, 11, 43, 20, 54, 5, 11, 24, 9, -20, 13, 5, 1, 26, 9, -25, -33, -79, -48, -45, -15, -8, -4, -23, -16, -43, -49, -10, 18, 15, 27, -5, 17, 9, 22, -6, -45, -26, -19, -15, 16, 1, 1, 12, 25, -11, 7, 8, -6, -1, -45, -13, 15, -46, 5, 19, 11, 48, 43, 37, 8, -7, 64, 37, -17, -23, -28, -5, -17, 12, 18, 29, 33, 58, 33, 46, 10, 8, -20, -8, 3, 12, 20, 28, 49, 78, 85, 106, 66, 38, 32, 21, -24, 5, 17, -18, -4, 5, -18, 8, -5, 23, 7, 15, 33, 20, 2, 51, 49, -4, -17, 19, 35, 11, 25, 24, 9, 2, 28, 8, -12, -5, 5, -4, -15, 19, -17, 20, -13, 14, -20, -12, -4, -6, 1, 0, -9, 3, 11, -5, 20, -20, -5, 13, 11, 13, -9, 8, 16, 13, -6, 5, 1, -1954, 2, -6, -16, -4, -19, 9, -14, 5, 37, 21, 22, 11, 25, 22, 1, 5, -1, 6, 7, -21, -12, -25, -24, -25, 2, -10, 2, -10, 4, 16, -9, -12, -55, -29, -31, -1, 5, -10, -31, -40, -8, 10, -63, 13, -43, -30, -4, -20, 7, -23, 28, 80, 22, -5, 15, 14, -6, -16, -24, 4, 66, 24, -25, -27, -53, -95, -91, -105, -77, -20, -11, -59, -64, -80, -21, 26, 6, -60, -34, 42, 36, -15, -3, 18, -2, 18, 14, 39, 40, 3, -47, -52, -30, -38, -45, -112, -25, -29, -30, -5, -36, 22, -48, -18, -16, 1, 8, -7, -55, -27, 2, 19, 12, 37, 9, 21, -1, -14, -66, -69, -42, 10, 78, -6, -2, -24, -2, -7, -45, -14, -41, -19, -18, 16, 42, -23, -31, -30, -14, -2, -2, 22, -11, 27, 23, -36, -64, -14, -4, 23, 18, -10, -10, 5, -51, -79, -95, -32, -71, -60, -48, -1, 59, -21, -28, -29, -4, -5, 13, -4, 30, 41, 30, -21, -58, -43, -33, -3, -28, -23, -5, -6, -53, -45, -18, -32, -46, -59, -34, -34, -9, -29, -58, -36, -10, 21, 27, 8, -4, 5, -20, -65, -88, -43, -5, -4, -26, -8, -2, -10, -25, 7, 30, -29, -74, -18, -32, -43, -26, -7, -67, -15, 20, 8, 33, 0, 12, 24, -24, -84, -87, -32, 8, 1, -40, -61, -44, -20, -14, 49, 16, -14, 0, -12, -29, -71, -115, -58, -29, -38, -31, 23, 2, 21, 22, -29, -26, -44, -7, 14, 50, -19, -47, -128, -71, 23, 61, 39, 9, 27, 21, -37, -91, -156, -130, -61, 2, -15, 6, -35, -73, 3, -27, 3, 46, 0, 44, 75, -11, -48, -105, -104, -18, 65, 48, 28, 8, 21, -29, -75, -115, -190, -99, -48, 8, 3, 8, -10, -74, -39, -57, -11, 0, -42, 19, 7, -76, -116, -110, -36, -11, 36, 31, 17, 45, 21, -26, -58, -122, -126, -89, -10, -24, 9, 2, 19, -39, -67, -48, -76, -34, -33, -21, -97, -154, -99, -18, 20, 21, 37, 50, 31, 34, -26, -30, -48, -107, -106, -75, 18, -25, 33, 6, -16, -33, -61, -53, -61, -52, -66, -33, -80, -102, -60, 16, 65, 44, 9, 10, 36, 8, -2, -47, -64, -93, -88, -80, 38, 32, 14, 3, -11, -39, -71, -69, -98, -54, -47, -17, -88, -104, -10, 59, 59, 57, 43, 40, 59, 38, 13, -63, -79, -130, -112, -75, 29, -3, -37, -21, 8, -19, -80, -98, -59, -64, -71, -32, -104, -94, 3, 13, 65, 39, 59, 46, 92, 24, 5, -48, -151, -156, -115, -82, 19, -1, 0, -7, 3, 1, -53, -101, -133, -124, -106, -97, -106, -75, 7, 2, 54, 67, 54, 91, 60, 20, -21, -132, -218, -181, -145, -49, -16, -40, 40, 6, -34, 19, -47, -83, -121, -140, -89, -73, -135, -34, -41, 3, 19, 58, 74, 81, 53, 26, -38, -133, -155, -144, -137, -70, -47, -30, -7, -10, -36, 31, -26, -115, -106, -100, -56, -97, -104, -49, -17, -6, -10, 34, 61, 55, 13, 6, -18, -136, -155, -133, -87, -61, -47, -51, -60, -20, -47, -33, -80, -94, -156, -72, -52, -107, -63, 0, -6, 1, -24, -10, 27, 28, 4, -23, -31, -84, -100, -99, -88, -56, -13, -52, -55, -58, -7, -7, -32, -137, -152, -44, -36, -50, 11, 4, -5, 10, -2, -8, 24, 13, 9, 4, -58, -129, -151, -158, -104, -96, -42, -46, -56, -46, -5, 38, -13, -98, -44, -41, -16, -5, -48, -21, 15, -4, -50, -27, -44, -72, -29, -28, -72, -140, -123, -116, -109, -120, -13, 6, -38, -28, -2, -44, -71, -97, -14, -7, 2, 1, -40, -40, -40, -64, -60, -42, -69, -77, -54, -68, -67, -109, -129, -55, -53, -46, 28, 32, 37, 12, 16, -56, -59, -140, -101, -62, -21, -5, 4, 16, -10, -20, -6, -35, -40, -16, -32, -36, -35, -55, -29, -20, -45, -68, -35, 37, 44, 6, 16, 3, -74, -58, -39, -31, -7, -14, 51, 35, -31, 12, -61, -94, -127, -97, -127, -139, -99, -87, -79, -32, -20, -24, -12, 23, 27, -14, -7, 2, -15, -33, -36, 30, 84, 128, 54, 30, -36, -25, 18, 40, 37, -20, -82, -60, -53, -52, -47, -11, 3, -9, -10, 20, 13, -9, 21, 4, 4, -12, 0, 16, -7, 18, 35, 23, 0, -48, -17, 29, 69, 4, 27, 11, 2, -16, -18, -10, -10, -12, 1, 6, 3, 20, 4, -3, 10, -9, -14, -1, -14, 10, 15, 4, -15, -16, 6, -17, -18, 15, -14, 7, 2, 9, 0, -2, 11, 4, 16, -18, 7, -16, -9, 322, 11, -19, 16, 12, -13, 31, 17, 42, 42, 16, 70, 29, -36, -10, 39, 13, -24, 39, 45, 42, 25, 26, 7, -5, -20, -20, -8, 4, -19, -16, -5, 12, -19, 24, -5, 6, 64, -16, -27, 38, 29, -1, 48, 9, -34, -30, -53, -21, -17, -37, -41, -54, -4, 18, -3, 12, 12, 5, -9, 16, -17, -11, 10, -3, -1, -28, -17, 10, 22, 22, -44, -34, -42, -73, -47, -28, -16, 0, 12, 31, 0, -2, -3, 10, -3, 32, 60, 50, 8, 65, 87, -38, 7, 23, -1, -27, 18, 23, 3, -34, -3, -34, -2, -13, -15, 7, 0, -21, -118, 10, 4, -16, 19, 44, 27, 53, 94, 82, 95, 26, 24, 20, -21, -27, 25, 18, 6, -2, -3, 1, 23, 16, -12, -5, -27, -50, -100, -33, 0, -14, 14, 53, 87, 105, 154, 128, 91, 46, 39, 27, -7, -27, -3, 17, 9, -6, -20, -12, 1, -17, -10, -18, -13, -65, -39, 36, -19, -21, -6, 53, 75, 73, 133, 113, 37, -3, 12, -1, -9, -16, 2, 29, 2, 25, -4, -12, -39, -45, -30, -76, -53, -83, -24, 16, -25, 14, -22, -6, 38, 75, 77, 64, 6, -9, -2, -21, -46, -17, 18, 30, 37, 75, 35, -2, -27, -17, -49, -69, -50, -61, 5, 31, -21, 17, 37, 34, -5, 47, 86, 27, 17, -35, -40, -55, -13, -42, 4, 36, 100, 106, 115, 62, 52, -2, -38, -61, -71, -33, -8, 10, 11, 10, 56, -10, 71, 119, 103, 45, -10, -28, -32, -22, -34, -14, 28, 21, 81, 149, 159, 153, 96, 40, 7, -47, -34, -39, -21, -22, 4, 29, 57, 43, 158, 118, 20, 10, -35, -35, 5, 9, -21, 0, 31, 31, 79, 114, 158, 167, 132, 116, 31, 6, -11, -23, -18, 10, -23, -3, 44, 106, 112, 105, 48, 26, -18, 0, 10, 14, 65, 14, 17, -27, -17, 4, 45, 111, 154, 151, 138, 88, 54, 8, 19, -6, -9, 17, 35, 102, 75, 73, 40, 18, -3, 44, 62, 14, 21, -10, -6, -52, -85, -72, -45, 58, 89, 143, 191, 183, 154, 56, 51, -25, -20, 2, 44, 107, 103, 136, 105, 47, 41, 57, 48, 48, -7, -45, -44, -78, -113, -74, -43, 35, 52, 84, 109, 170, 169, 138, 125, 76, -20, -19, 38, 82, 116, 168, 127, 99, 49, 14, 22, 13, -1, -45, -62, -108, -118, -76, -42, 23, 0, 12, 30, 87, 174, 127, 128, 100, 17, 12, 33, 46, 56, 105, 67, 92, 20, -14, -8, -39, -26, -37, -50, -108, -108, -29, -14, 34, 10, 1, 25, 58, 138, 140, 114, 61, 49, 23, 23, -86, -71, -32, 24, 47, 11, -27, -23, -7, -15, -22, -51, -109, -55, -6, 28, 36, -4, -25, -7, 60, 110, 93, 42, 76, 63, 37, -1, -44, -48, -49, -24, 23, -9, -45, -35, 5, 27, 75, -15, -44, -22, 6, 31, -5, -36, -63, -15, 12, 113, 31, 18, 91, 14, 22, 5, -73, -101, -36, 23, 13, -15, -34, 23, 43, 55, 67, 39, -4, 22, 0, -20, 5, -33, -29, -25, -36, 67, 46, 13, 6, 31, 16, -24, -64, -100, -7, 48, 24, -12, 4, 8, 50, 60, 13, -6, -5, -28, -10, -16, -2, -13, -17, 21, -5, 14, 48, -7, 35, 50, -12, -15, 10, -84, 3, 47, 46, 39, -12, 3, 47, 7, 6, -11, -33, 12, 9, -2, 11, -3, 33, 36, 32, -5, 29, 41, 16, 26, -18, 8, -47, -60, -8, 13, 43, 42, 16, -18, 2, -13, -6, -6, -28, -27, -37, -5, -8, 29, -4, -31, 3, -11, 27, 28, 14, -10, -1, 20, -68, -27, 42, 51, 25, 23, 3, -15, 36, -9, -6, -4, -29, -42, -49, -28, 1, 35, 26, -21, -16, 12, 26, -9, 14, 4, -15, -33, -45, -51, -35, 29, 28, 6, 4, -4, 7, -14, -45, -49, -49, -21, -34, -9, 7, 21, 5, 26, 14, -3, -16, -29, 37, -14, 16, -19, 20, -3, -24, -32, -13, -15, 13, 15, -26, 11, -27, -43, -8, 31, 8, 82, 104, 94, 26, 14, 4, -15, -12, -10, 25, -19, -20, -9, -5, 19, 32, -4, 13, 24, -1, -19, -49, -36, -27, -31, 42, 22, 47, 56, 57, 58, 38, 5, 0, 18, -25, 12, 6, -10, 7, -11, -15, 13, 16, -3, 8, -23, -4, -12, -28, 42, 17, -6, -27, 10, -27, 14, 17, 10, 7, 18, 10, -12, -1, 17, 16, 2, -14, -3, 17, -18, 17, 17, 14, -12, 9, 18, -2, -15, 20, 4, -7, 8, -14, -5, 0, 8, -5, -13, 18, -8, 10, -20, 1, -20, -8, -1311, -20, 9, 0, 15, 2, -10, -27, -9, -34, -25, 18, 26, 24, -30, 31, 9, 48, 25, 29, 18, 14, -1, 16, -14, 19, 21, 2, -15, 2, 0, -4, 9, -23, -54, -88, -100, -40, -49, -76, -61, -18, -13, -36, -24, -13, 13, 21, -2, -27, -74, -76, -85, -17, -19, -14, 19, 14, 26, 30, -17, -29, -103, -52, -52, -61, -74, -26, 46, 27, -13, -50, -8, 16, -8, -4, 10, 33, 3, -35, -2, 29, -40, 10, 12, 5, 43, 48, 68, -20, -2, -34, -23, -16, -25, 0, -34, -47, -8, -19, 0, -16, -15, -20, 12, -18, -36, -39, 4, -46, -1, -5, 5, -18, 15, 7, -1, -41, 31, 40, 28, -12, -22, -29, 4, -19, 0, 34, 30, 38, 14, 20, 12, -11, 1, 9, -1, -60, -31, 12, -4, 3, -3, 6, -15, 9, 16, 41, 8, 14, 36, -13, 18, -23, 21, 27, 3, -13, 9, 7, 12, -10, -23, 25, 31, 7, 30, 9, 11, -21, 36, 4, -5, 35, 9, 16, -9, 27, 24, 14, -16, -10, 14, 25, 39, 3, -21, 16, -23, -38, -12, 27, -12, 20, 18, 16, -18, -6, 46, 3, -51, -22, 5, 10, -19, -14, -10, -11, -13, -18, 16, 5, 3, 14, -8, -19, -10, 0, 8, 13, 46, 25, -15, -23, 16, 35, 34, 28, -20, -30, 4, -20, -38, -16, 10, -33, -21, -32, -7, 37, 52, 47, 2, -4, 17, 2, 6, -18, 23, 28, -18, -22, -5, 61, 17, 56, 11, 39, 4, -37, -18, 3, 25, 4, -12, -58, -13, 35, 52, 29, 13, 1, 15, 16, -4, -1, 26, 21, -24, 10, 20, 72, 44, 48, 26, -4, 6, 10, -2, 1, -6, -43, -52, -32, 16, 55, 67, 64, 62, 68, 33, 4, 56, 14, -2, -11, -11, -32, 14, 60, 67, 44, 42, 45, -4, 48, -5, 17, -11, -35, -29, -12, -9, 42, 39, 62, 83, 80, 44, 54, 38, -1, -70, -20, 6, -30, -18, 62, 40, 52, 65, 25, 14, 31, -26, -10, -22, -31, -5, -8, 25, 79, 74, 114, 101, 41, 23, 10, -24, -89, -102, -38, -35, -25, 18, 49, 90, 59, 32, 37, -1, 22, 2, -12, -11, -39, -44, -10, 6, 78, 84, 72, 50, -11, -95, -147, -185, -208, -179, -90, -6, -12, 23, 31, 60, 68, 82, 4, -7, -2, -9, 5, -45, -41, -37, -32, 15, 28, 29, -58, -121, -210, -296, -345, -271, -237, -176, -100, 10, -13, 11, 29, -29, 65, -5, -52, -23, 5, -12, -51, -74, -82, -36, -28, -60, -79, -125, -232, -305, -315, -253, -219, -146, -98, -92, -82, -26, -3, -9, -24, -89, 1, -39, -47, 3, 20, -42, -42, -47, -70, -17, -57, -105, -174, -179, -133, -152, -103, -36, -53, -24, -20, -53, -91, -15, 11, -4, 15, 16, -45, -77, -25, -4, -24, -61, -69, -35, 1, -39, -44, -76, -92, -83, -47, 22, 31, 44, 43, 40, 44, -48, -80, 26, -1, 21, 14, -5, -100, -139, -13, 2, -12, -65, -31, -27, -18, -18, -2, -5, -7, 11, 11, 27, 69, 49, 28, 11, 62, 9, -15, 30, 16, 24, -15, -50, -131, -139, 1, 7, -37, -15, -3, -41, -5, -28, -3, 58, 36, 29, 37, 72, 32, 41, 17, 21, 45, 47, -2, 13, 53, -10, 33, -7, -91, -67, -34, 0, -17, 19, 28, -4, -7, -23, 10, 34, 46, 35, 27, 45, 24, 36, 40, 30, 23, 19, 15, -8, 34, -18, 10, 8, -46, -66, -30, -26, -12, -3, -17, -10, -8, -1, -20, 11, 3, -28, 3, 21, 4, -10, 7, 13, -39, -5, -31, -25, 37, -13, 7, 11, -9, -14, 6, -22, -15, -27, -57, -30, -44, 5, -3, -41, -15, -27, -9, 2, -17, -2, -11, -7, 9, 4, 5, 41, 1, -11, 11, -14, -5, -36, -21, 1, -19, -2, 20, -6, -35, -21, -59, -38, -48, -31, -32, -8, -14, -33, -19, 33, -21, -11, -21, 27, -4, 1, 12, 16, -7, 45, 18, 32, 47, 28, 27, -28, -8, 15, -36, -27, -4, -1, -5, 5, 53, -2, 9, 45, 14, -10, 15, 21, 7, -17, 10, 16, 54, 61, 35, 32, 58, 44, 39, 51, 27, 66, 37, 37, 31, 63, 50, 76, 88, 77, 4, 27, 22, 12, -11, 6, -1, 17, 19, 5, 0, 9, 34, 21, 25, 32, 5, -14, 21, 33, -11, -6, -27, -1, -15, -27, -7, 14, 0, 12, 19, -2, 12, -10, -12, -16, 4, 1, -6, 8, -2, -7, -17, 13, -16, -6, 18, -2, -6, 19, 7, 14, -4, 13, 6, 2, 7, -2, -9, -15, -1, -12, -16, 17, -1131, -2, 2, -8, 20, 15, 31, 34, 51, 49, 73, 91, 62, 26, 36, 77, 20, 6, 18, 47, 5, 16, -15, 8, 25, -5, -20, -3, -9, 7, -14, -2, -9, -56, 25, 15, -21, 34, 0, 0, 9, 46, 29, -17, -27, -40, -10, 79, 89, 83, 43, 32, -7, -8, 9, 17, -19, -6, -17, 27, -35, -16, -31, -43, -3, -14, 2, 22, 2, -34, 6, -68, -43, -45, -58, -14, -16, 14, 16, 32, 67, 42, -5, 20, 3, -15, 20, -8, -39, 15, -29, -15, 3, 11, 4, 17, -6, -6, -7, -29, -59, -24, -13, -66, -42, 18, 36, 58, 5, -43, 16, -14, -3, -4, 14, -7, -22, -34, -40, -64, -69, -38, 6, 52, 18, 19, 28, 12, -11, -23, -3, -19, -33, 19, 8, -8, -60, -84, -43, 11, -3, -6, 24, -38, -25, -57, -63, -65, -84, -48, -50, 30, 15, 37, 18, -18, -23, -19, 4, -1, 24, 0, -35, -33, -88, -87, -42, -10, 8, 15, -21, -29, -27, -68, -102, -59, -114, -90, -91, -48, 1, -31, -29, -49, 3, -5, 17, -5, 14, -60, -98, -90, -95, -127, -68, -7, 9, -4, -13, -24, -41, -136, -122, -83, -143, -162, -116, -43, -34, -47, -43, -17, -22, 10, -12, -46, -18, -63, -135, -135, -98, -140, -34, -38, 2, 21, -8, -28, -123, -179, -157, -116, -125, -143, -130, -87, -104, -84, -25, -28, -18, -38, -68, -93, -103, -122, -130, -115, -11, -21, -23, 45, 6, 16, 43, -26, -113, -143, -93, -37, -103, -100, -82, -77, -90, -60, -15, -22, 5, -51, -96, -146, -174, -151, -132, -85, 11, -28, 5, -9, 19, -59, -10, -22, -61, -59, -11, -16, -28, -43, -27, -12, -41, -25, 1, 49, -1, -72, -76, -97, -30, -40, -78, -45, 4, -25, -34, 22, -19, -61, -86, -91, -63, 0, -9, 16, 25, 9, 4, 38, 45, 45, 65, 24, -6, -62, -56, -33, 10, 25, 3, -15, 72, -1, -29, -3, -1, -19, -32, -53, -78, 33, 68, 39, 31, 41, 54, 82, 71, 40, 34, 39, -15, -37, -17, 3, 15, 8, -14, 20, 66, 38, 47, 28, -34, 6, -65, -22, -58, -9, 40, 60, 81, 78, 60, 30, 68, 62, 49, 9, 0, -3, 16, 11, 33, 37, 22, 48, 92, 114, 92, 51, -23, -23, -46, 2, -70, -35, 54, 63, 26, 17, 11, 18, 56, 75, 27, -34, -34, -27, 36, 9, 3, 21, 5, 25, 114, 75, 91, 59, 7, 42, -41, -62, -94, -26, 38, 13, 16, 16, 27, 29, 85, 77, 14, -46, -15, -16, 18, 23, 38, 35, -22, -1, 48, 60, 70, 53, 38, 72, -65, -63, -80, -74, 18, 31, -21, -6, -45, 21, 48, 74, 27, -27, 17, -3, 22, 7, 50, 38, -5, 12, 7, 49, 91, 9, 41, 34, -38, 5, -34, -15, 1, 10, -6, -20, -16, -13, 29, 69, 40, 8, -15, -6, -20, 26, 35, -2, -8, 25, 1, 23, 18, 61, -11, 17, -14, -30, -7, -19, 30, 28, -6, -24, -7, 3, 13, 51, 47, 0, -13, -7, -6, 14, 30, 15, 11, 33, -6, 12, 23, 66, -12, -12, 39, 19, -5, 42, 40, -8, 11, -27, 1, -11, -40, -4, 10, -25, 3, -1, -4, 35, 62, 2, 4, 28, 43, 53, 48, 37, -22, -28, 52, 16, 49, 47, 27, 7, 28, 15, 7, 36, 8, -10, -8, 6, -9, 3, -11, 34, 13, 16, 18, -5, 11, 95, 69, 2, 14, -3, 33, -32, 2, 26, 5, 39, -9, -53, -7, 22, -13, -9, -13, -26, 11, 9, -20, 10, 18, -1, 7, 45, -16, 44, 3, -32, 11, -19, -66, -52, -1, 21, -33, -53, -107, -66, -60, -77, -60, -6, -49, -54, -16, -49, -79, -38, -18, -43, -45, 25, -45, 12, 21, 19, 2, -27, -44, -52, -23, 1, -7, -18, -10, -26, -88, -90, -82, -111, -149, -142, -92, -116, -143, -123, -125, -107, -68, -26, -46, 39, 9, 16, -5, -5, -3, -19, 22, -11, -48, -45, -80, -60, -56, -79, -128, -177, -206, -202, -168, -166, -114, -124, -141, -115, -40, -40, -31, -15, 18, 9, 20, -17, -1, -19, -6, -61, -73, -59, -66, -76, -68, -55, -120, -124, -127, -122, -95, -108, -73, -81, -27, -35, -39, -14, -34, -9, -2, 10, 6, -19, 9, 20, -8, -50, -59, -29, -59, -54, -38, -60, -59, -65, -26, -63, -59, -35, -34, -34, -20, -21, -36, -25, 14, -17, -11, 14, 7, 14, -15, 4, 12, -10, 5, 20, 9, 2, 8, -17, 4, -16, 19, -21, 5, -21, -21, -5, 7, 2, -14, -17, 10, 16, 4, 3, -5, -1159, -10, 12, -11, 21, -20, -62, -49, -81, -67, -56, -62, -87, -75, -112, -86, -76, -60, -52, -53, -51, -27, -27, -1, 8, 0, 6, -17, -11, -12, -10, 3, -29, -31, -108, -138, -105, -91, -125, -126, -105, -110, -181, -177, -167, -108, -145, -123, -108, -123, -92, -47, -48, 3, 9, 13, 0, 16, 30, 23, -42, -50, -91, -84, -23, -47, -62, -74, -105, -93, -120, -194, -221, -197, -233, -185, -138, -165, -81, -64, -27, -16, -4, -7, -12, -14, 6, 24, 29, -52, -39, 22, -11, 10, 28, -32, -60, -62, -101, -124, -95, -88, -61, 7, -4, -6, -12, -6, 0, 1, 14, -20, 11, 13, -5, -30, -41, -88, -12, 59, 25, 28, 16, -35, -75, -46, -29, -67, -33, 8, 29, 39, 55, 57, 35, -10, -19, 42, 71, -8, -7, -10, 15, -42, -43, -18, 20, 58, 0, 2, 6, -22, -14, -26, -56, -52, -19, 6, 3, -15, -26, -23, -25, 9, -12, 65, 70, 3, 10, -12, 58, -29, -56, -22, 30, 4, -8, 27, 29, 22, -3, -10, -28, 1, 25, 9, -7, 15, -4, -38, -50, -24, 20, 129, 70, 7, 2, 8, 21, -35, -48, -40, -13, 44, 21, 2, 69, 19, 38, 53, 46, 32, 46, 66, 7, 34, 30, -6, -18, 7, 84, 141, 35, 25, -1, 27, 9, 25, -51, -43, 8, 9, -19, -15, 46, 21, 62, 76, 45, 27, 20, 35, 5, 26, 6, 31, -4, 32, 61, 82, -10, -43, 10, 63, -38, 40, 27, 14, 42, 52, 4, -21, 46, 37, 51, 54, 4, 9, 3, 0, 10, 1, 21, 11, -1, -11, 15, 52, 14, 18, -22, 64, 46, 77, -11, 18, 83, 47, 25, 13, 32, 39, 21, 12, -31, -28, 12, 27, 50, 29, 26, 26, -10, 6, 0, 10, 50, 14, 17, 59, 132, 135, 50, 72, 51, 61, 65, 43, 16, 11, 44, 28, -42, -39, 7, 48, 6, 44, 28, 32, -3, 33, 19, 45, 60, 9, 16, 37, 106, 78, 75, 42, 33, 32, 33, 2, -21, -6, -18, -58, -65, -25, 24, 15, 27, 42, 40, 40, -3, 42, 16, 34, 45, 16, 15, 27, 25, 23, 65, 44, 23, 9, 0, -9, -21, -11, -45, -60, -79, -22, 7, 14, 41, 39, 35, 35, 9, 19, 1, 20, -21, 9, 6, 4, 7, -9, 5, 38, 9, -24, -59, -21, -5, -32, -34, -52, -95, -44, -8, -9, 4, 27, 28, 21, 0, -53, -84, -4, -37, 7, 10, -39, -53, -70, -29, -51, -15, -56, -78, -74, -23, -43, 1, -33, -70, -8, 30, -28, -37, -31, -34, -29, -48, -42, -77, -30, -17, -18, 6, -33, -93, -136, -140, -98, -100, -78, -88, -39, -36, -6, 12, 11, -44, -29, -31, -66, -47, -41, -23, -40, -39, -33, -34, 5, -20, 15, 14, -24, -69, -146, -137, -115, -65, -66, -64, -36, -47, 43, 67, 60, 0, -28, -67, -86, -70, -79, -35, -43, -43, -1, 32, 37, -26, -48, -8, -63, -79, -153, -165, -130, -80, -52, -6, -19, -28, 6, 79, 53, -10, -22, -49, -101, -69, -62, -46, -32, -24, 24, 25, 6, -18, -66, -5, -46, -76, -217, -164, -77, -67, -22, -3, -33, 6, 24, 51, 48, 15, -32, -52, -91, -76, -58, -42, -28, -3, 32, 45, 59, 17, -25, 31, 19, -23, -99, -54, -23, 16, -18, -1, -18, -12, 12, 12, 8, 12, -40, -88, -85, -108, -83, -66, -43, 2, 48, 52, 16, 16, 13, -17, 0, -18, -55, -1, 7, -18, -21, -43, -38, -32, 4, 14, 10, -13, -35, -104, -105, -108, -87, -64, -32, -18, 31, 90, 39, 31, 38, 16, 24, 13, -38, -5, 30, -28, -25, -48, -29, 35, 24, 54, 24, 48, -1, -54, -33, -15, -63, -42, -44, 8, 5, 63, 9, -17, -13, 2, 17, -35, -82, -98, -63, -29, -35, -18, -26, -17, 7, 28, 34, 21, 35, -7, 8, 54, 49, 63, 59, 48, 52, 7, -64, -34, -21, -11, 5, 0, -46, -43, -89, -69, -45, -58, -49, -54, 32, 64, 39, 62, 34, 66, 97, 81, 72, 88, 65, 26, 29, -15, 46, -27, -1, 21, 14, -5, -33, -11, 14, -20, -2, -17, -35, -37, -7, -44, -47, 44, 55, 80, 85, 69, 17, 10, 14, -29, -7, 39, 21, 5, -17, 9, 8, 2, -4, 1, 27, 24, 2, -11, -26, -22, 12, -15, -24, -2, 8, 25, 0, -13, -38, -32, -10, -22, 3, 2, -11, 5, 14, 6, 6, -9, -1, -14, -11, 2, 16, -3, 9, 11, 15, -18, 12, 8, -4, -15, -6, 9, -8, -1, 4, -1, -20, 4, 17, -11, -8, -9, -1842, -2, 12, 10, -2, 8, -3, 2, 11, 5, 2, -3, 45, -8, -52, 23, 0, 45, 37, 14, -26, -15, 21, 8, 14, 0, 17, 5, 1, 17, -13, -7, -21, -53, -12, -51, -87, -111, -108, -111, -78, -22, -32, -65, -68, -51, -27, 45, 69, 43, -44, -55, -90, 8, -6, -3, -17, -5, 18, 32, -21, -37, -69, -82, -176, -180, -148, -118, -77, -71, -46, -61, -43, -28, -76, -4, 3, 7, -36, -6, 47, 64, -43, -17, 16, -4, 30, 65, 20, -71, -50, -74, -105, -111, -129, -73, -107, -46, -17, -31, -15, -28, -44, -54, -50, -48, -2, 13, 2, -95, -5, -7, 14, 0, 40, -29, -60, -79, -41, -29, -38, -69, -67, -46, -14, -23, -37, 3, -11, -47, -65, -39, -93, -33, 9, 74, -7, -65, -24, 10, -14, -11, -6, -46, -47, -63, -23, 4, 1, 23, 4, -14, -4, -18, -27, -54, -51, -56, -26, 5, 1, -10, 44, 84, 54, 3, 28, 3, 7, 13, 17, 9, 36, 11, -18, 6, 30, 22, 7, -2, -8, 7, 26, -31, -6, -23, 0, -28, -33, -4, 34, 57, 11, 1, 16, -7, 19, -10, 67, 18, 23, -9, -14, -4, -19, 21, 36, 22, 28, 7, 59, -20, 36, 8, 24, -17, -7, -8, -10, -31, 22, 34, 20, -39, 21, 38, 72, 96, 19, 6, -2, -1, 14, -24, -22, 18, 4, 20, 51, 40, 82, 43, 1, 29, -24, 25, -26, -33, -3, 17, 6, -25, -2, 29, 86, 183, 67, 27, 15, 22, -19, -26, 20, -11, -26, 22, 68, 82, 81, 22, 1, -3, 25, -12, -52, -30, -21, 22, -57, 4, 23, 23, 85, 180, 72, 34, 19, -8, -19, -79, -31, -43, -12, 28, 54, 81, 60, 42, 17, 1, -10, -23, 0, -40, -76, -52, -52, -8, -3, 59, 39, 91, 33, -21, -29, -16, -37, -56, -51, -18, -5, 29, 70, 84, 84, 58, 22, 30, 20, 12, 11, -26, -83, -68, -18, -25, -10, 11, 35, 55, 11, 59, 38, 0, -41, -53, -42, 3, 5, 47, 41, 51, 40, 35, 0, -30, -30, -33, -71, -72, -112, -69, -31, -3, 9, -1, 36, 49, 46, 81, 59, -18, -25, -7, -30, -2, 23, 25, 39, 5, 27, -4, -32, -109, -97, -73, -73, -77, -113, -54, -1, -3, 2, -10, 21, 87, 78, 62, -4, -17, -37, -40, -10, 15, 7, 11, 1, -5, -46, -97, -161, -149, -145, -115, -78, -101, -90, -44, 28, -3, -10, 41, -14, 37, 24, 16, -15, -27, -47, -45, -23, -19, -10, 20, 20, -68, -75, -147, -163, -119, -35, -69, -99, -130, -60, -73, 8, 25, 13, -24, -104, -51, -70, -21, -18, 10, -38, -79, -42, -24, 9, 41, 2, -79, -93, -85, -56, -27, 6, -55, -53, -78, -101, -94, 14, -1, 19, 13, -31, -59, -59, -57, -51, -18, -62, -67, -42, 28, 16, 50, -15, -59, -89, -50, -35, 19, 2, -18, -40, -34, -56, -79, 21, 36, 13, 10, -48, -137, -93, -61, -16, -14, -50, -43, -19, 1, 10, 27, 1, -18, -40, -14, 12, 20, 14, 25, -19, -4, -17, -46, 8, 51, 25, -33, -59, -158, -103, -46, -9, -11, 17, -17, 18, 11, -43, -1, -4, -34, -5, 17, 62, 58, 25, 35, 1, 41, 63, -27, -16, 44, -6, 10, 5, -121, -57, -17, -3, 12, 51, 23, 0, -16, -46, -45, -49, -6, 9, 47, 50, 12, 32, 37, 24, 6, 66, 17, 25, 32, -7, 7, -3, -35, -46, -41, -25, -24, -10, -11, 0, -31, -36, -57, -62, -21, 39, 57, 65, 15, 18, 51, 76, 50, 29, 2, -13, 2, 0, 11, -15, -57, 6, -27, -65, -35, -81, -80, -80, -70, -22, 3, -3, 7, 21, -12, 13, 9, 46, 5, 47, 61, 50, -38, 62, 8, 10, -23, -69, -71, -30, -58, -40, -34, -53, -35, -60, -43, -29, 9, 20, 28, -19, -18, -20, -22, -24, 11, 29, 25, 38, -7, 15, -12, -3, 8, 5, 6, 38, 22, -6, 12, -22, -1, -46, -11, 26, -2, -30, -7, -44, -62, -10, 21, -14, -5, 40, 2, 36, -2, 8, -8, 1, -19, -13, 52, 48, 46, 48, 64, 32, 42, -18, 60, 88, 144, 135, 102, 75, 118, 97, 93, 87, 56, 81, 34, 21, 18, 23, -13, 18, -1, -1, -10, 10, 34, 55, 65, 80, 61, 68, 12, 21, 51, 1, 50, 78, 65, 64, 33, 53, 36, 25, -11, 6, -18, -7, 3, -14, -19, -18, -16, -5, 18, 1, 3, -20, -9, -1, 4, 2, -14, -14, 24, 30, -13, -21, -15, -8, -17, 20, -16, -16, 2, -4, -7, 7, -64, 8, -18, 11, -17, -43, 8, -5, 10, 47, 41, -13, 5, 54, 106, 41, 73, 28, 50, 62, 24, 11, 24, -16, 3, -20, -1, 13, -15, 5, -15, -14, 14, 37, 58, 61, 131, 107, 122, 121, 137, 131, 174, 172, 153, 130, 111, 124, 113, 112, 87, 43, 86, 16, -1, -5, -2, 19, -23, 0, 38, 61, 41, 53, 91, 121, 92, 67, 46, 47, 57, 58, 81, 78, 68, 80, 115, 88, 73, 77, 69, 4, 39, 15, 4, 13, -31, -56, -4, 60, 25, -11, 27, -6, -6, 10, 24, 15, 9, 52, 41, -25, 39, -5, 54, 67, 86, 116, 129, 95, 4, -7, -10, -19, -35, 2, 61, 47, -9, -75, -35, -57, -42, -2, -13, 19, -27, -8, -40, -35, 0, -18, 14, 11, 35, 53, 41, 62, -16, 4, -3, 31, -13, 14, 45, -9, -74, -124, -81, -75, -56, -47, -27, -34, -46, -51, -51, -39, -55, -59, -31, -9, 22, -28, -6, 19, -23, -17, -10, -13, -7, 7, 24, -45, -84, -99, -25, -45, -12, -42, -23, -54, -94, -51, -36, -49, -56, -64, -20, -10, 29, 3, -12, -5, -17, -32, -1, 21, -80, 30, 19, -28, -47, -55, -50, 33, 6, 22, -25, -32, -38, 1, -16, -32, -35, -62, -7, -46, 5, 28, -11, -16, 20, 16, -18, -27, -85, -19, -18, -40, -32, -25, 11, 37, 41, 7, -19, -25, -16, 8, 21, 2, -33, -8, 16, 8, -13, 6, 15, -47, 75, 9, 6, -57, 5, -55, -53, -53, 25, -55, -35, 19, 27, 48, 9, 4, -43, -43, -15, 35, 25, -7, 10, 30, 6, -4, -2, -56, 36, -14, 38, 17, -43, -89, 13, -18, -17, -28, -11, 7, 17, 52, 16, -19, -41, -58, -24, -6, 4, 9, -1, 0, -10, 31, 43, -21, 9, 23, 12, -10, -112, -81, 7, 1, 3, -52, -7, -26, 20, 12, -4, -51, -83, -93, -36, -4, 22, 15, 23, 2, 33, 28, 57, 0, 2, 27, -17, -52, -80, -40, 29, -2, -13, -29, 8, -23, 19, -16, -40, -81, -113, -74, -41, -16, 3, 26, 17, 10, 21, 74, 25, -17, -39, 3, 4, -16, -59, -48, 5, -7, -8, 18, 9, -16, -9, -4, -83, -55, -48, -43, -18, -3, -3, 23, 7, 45, 17, 67, 54, 22, -60, -26, -28, -43, -57, -32, -40, -37, -11, -35, -8, -11, -35, -23, -76, -61, -22, 23, 6, -4, 16, -4, 10, 18, 34, 72, 135, 29, -59, -31, -1, -46, 51, -42, -29, 37, -2, 8, 5, 30, -8, 5, -41, -10, -7, 16, -41, -19, 3, -1, -11, -30, 21, 34, 69, 32, -42, -61, -10, 10, 73, 46, 83, 32, 46, 42, 55, -20, 16, 58, -11, -14, 11, 19, 0, -4, -32, -9, -1, -20, 25, -20, -3, -12, -37, -19, 0, -12, 29, 58, 54, 48, 41, 42, 14, 2, 39, 45, 55, 33, 54, 6, -23, 0, 7, -4, -20, -13, -28, -45, -41, 4, -5, -63, -11, -22, 20, 54, 74, 2, 10, 16, 16, 16, 71, 66, 75, 64, 62, 19, 27, 28, -6, 4, -10, -17, -48, -85, -99, 14, -10, -15, -38, 8, -16, -52, 0, 12, -1, 27, 37, 25, 97, 92, 107, 70, 46, 54, 50, 40, -2, 6, -16, -43, -81, -102, -59, -34, -29, 5, 9, -2, -42, -9, -16, -7, -18, 30, 21, 43, 67, 58, 74, 85, 56, 52, 81, 45, 19, -11, -24, -88, -69, -73, -73, -32, 0, -52, -1, 12, 35, -18, -24, -12, 14, 31, 33, 37, 20, 19, 9, 29, 32, 64, 38, 40, 1, -49, -91, -84, -49, -15, 2, 33, 13, -7, 16, -18, 13, -12, -40, -67, -29, -16, -18, -48, -71, -55, -80, -55, -27, 34, 5, 2, -61, -108, -141, -58, -25, 6, -22, 4, -41, -20, 6, -10, 58, -3, 0, -21, -43, -50, -82, -48, -54, -57, -66, -14, -3, -21, -9, -18, -63, -78, -83, -76, -74, -38, -4, 47, 10, 15, 12, -19, 16, 17, -47, -54, -76, -53, -22, -81, -70, -34, -27, -33, -19, -50, -8, -16, -62, 0, 2, -17, -21, 0, 26, 19, 11, 16, -2, -12, 9, -13, -69, -41, -103, -74, -80, -31, -44, -98, -47, -142, -94, -77, -34, -44, -87, -61, -42, 14, -41, -16, 29, 32, 6, 2, 2, 6, -12, -1, -15, 0, -2, -1, -45, -16, -54, 30, 21, -2, -16, 2, 17, 3, -43, 10, -12, -22, 11, 8, 17, -7, -18, 13, 14, -17, 6, -5, 1, 13, 0, 11, 15, -17, 20, 4, -16, 17, -1, -21, 15, 7, 19, 1, -3, 2, -18, -3, 7, -11, -8, -18, 1, -717, 1, 8, 17, -20, 34, 35, 30, 71, 53, 50, 115, 113, 59, 104, 64, 30, 30, 63, 49, 47, 17, 35, -5, -10, 1, 1, -18, 0, 13, -13, 21, 21, 33, 108, 72, 114, 114, 111, 109, 86, 97, 195, 122, 64, 120, 145, 143, 116, 140, 124, 93, 53, 18, 6, 7, 11, 13, -34, -1, 37, 61, 50, 96, 86, 97, 57, 54, 8, 2, 30, 43, 83, 59, 53, 105, 129, 95, 55, 104, 43, 1, 16, 4, 7, -20, -29, -23, -7, 56, 29, 33, 41, -16, -45, -6, -19, -35, -19, 9, -12, -18, 33, 2, 29, 44, 76, 73, 84, 35, 15, -4, -10, 10, 4, 27, 58, 25, -7, -24, -33, -88, -61, -45, -24, -23, -43, -32, -33, -40, -34, -43, -5, 36, 6, 53, 49, -12, -15, -14, -13, 4, -17, -6, 13, -4, -14, -75, -53, -76, -59, -20, -26, -29, -6, -26, -47, -93, -44, -36, -46, 9, -31, 1, -11, -42, -57, 15, -6, -2, -62, 29, 4, -31, -43, -55, -26, -64, -32, -38, -27, 4, -22, -39, -51, -89, -38, -56, -53, -17, -21, -78, -86, -29, -2, -26, -13, 27, -27, 12, -45, -46, -56, -114, -51, -8, -33, -17, -14, -28, 0, -18, -52, -41, -60, -94, -90, -84, -73, -82, -92, -91, -25, 32, -3, 39, -20, -26, -99, -137, -107, -70, -28, 29, 15, 9, -20, -38, -16, 18, -14, -9, -23, -37, -61, -88, -93, -100, -94, -42, 72, 61, -16, -12, 51, -81, -206, -180, -126, -42, -2, 29, 20, 14, -6, -6, 14, 63, 44, 37, 56, 23, -3, -49, -75, -55, -81, -28, 51, 19, 60, -23, -53, -120, -103, -149, -61, -44, 12, 53, 61, 37, -14, 8, 16, 41, 51, 71, 69, 89, 77, 39, 27, 11, -21, 20, -12, 37, 20, -45, -84, -201, -118, -103, -59, -13, -6, 42, 54, -8, -31, -35, 8, 17, -4, 16, 40, 76, 69, 58, 39, 30, 1, -31, 26, 43, 10, -48, -98, -129, -119, -87, -73, -4, 39, 48, 77, 0, -45, -45, -29, -30, -33, -32, -31, 14, 58, 57, 97, 67, 36, -29, -26, 34, 3, -50, -100, -59, -87, -97, -74, -6, 30, 26, 38, -7, -47, 4, 0, -26, -89, -114, -35, -5, -2, 11, 38, 37, 51, 26, 42, 14, -22, -31, -46, -26, -78, -74, -55, 5, 21, 23, 23, 4, -6, 19, 5, -34, -142, -157, -88, -37, -5, 54, 29, 43, 103, 39, 41, -13, 4, 4, -8, -15, -73, 63, 38, 14, 59, 62, 62, 66, 39, 68, 61, -54, -113, -69, -56, -30, 15, 27, 24, 56, 67, 56, 36, -2, 3, 56, 50, -20, 27, 36, 70, 81, 92, 36, 64, 76, 39, 69, 56, -3, -75, -37, -25, -28, 27, 17, 36, 23, 12, -3, 44, 1, 34, 30, 12, 20, -36, -24, 14, 27, 63, 60, 28, 23, 16, 24, 19, -18, -57, -48, -67, -57, -11, 10, 16, -10, -26, -19, 60, 69, 5, 22, 2, -65, -77, -76, -7, 12, 6, 27, 23, 27, 23, 21, -5, -7, -54, -49, -49, -22, -1, 0, 36, -19, 18, 4, 39, 71, 4, -6, -54, -160, -80, -43, 14, 18, 29, 18, 36, 31, 29, 11, 1, 25, -4, -38, -48, 4, 36, 19, -47, -58, -13, 41, 20, 5, -40, -30, -80, -143, -91, -5, -29, -7, 66, 65, 49, 31, 31, 21, 25, 10, -11, -24, -9, -18, -16, 5, -12, -59, -35, 24, 27, 37, 5, -13, -28, -62, -21, -17, -31, 15, 41, 33, 30, 14, -6, 4, 15, 23, -15, -9, 4, -14, -18, -6, 26, 9, 21, 40, 68, -12, -9, -22, -14, -73, 22, 9, 10, 4, 5, 11, -15, -62, -100, -53, -10, -12, -20, -63, -80, -30, -17, 40, 36, 33, -6, 20, 46, -2, -5, -39, 4, -15, 33, 65, 75, 29, 43, 66, 39, 11, -2, -19, -29, -57, -88, -114, -164, -175, -98, -10, -1, 39, 45, 80, 41, -16, 11, 9, -10, -6, 10, 0, -20, -24, 8, 36, 62, 11, 6, 6, -57, -17, 7, -65, -47, -25, 21, 50, 8, -24, 48, 62, 32, -3, 8, 1, 15, 16, 7, -2, 31, 4, 5, -18, -9, -23, -6, -17, 4, -11, -31, -8, -18, 28, 69, 26, 39, 14, 45, 28, 3, 14, 13, 18, -9, 16, -5, 35, 43, 50, 75, 37, 36, -10, -34, 32, -7, 36, 20, 36, 54, 42, 29, 36, 23, -9, 12, 20, -16, 8, -18, -11, 10, -6, 14, -3, -1, -13, 0, 7, -5, -2, -9, 9, 5, -7, 11, -10, -15, 2, -7, -18, -9, -19, -5, -14, 19, 0, 6, 1510, -17, 14, 8, -12, 22, 16, 36, 51, 32, 27, 24, 6, 3, 11, 72, 67, 58, 65, 26, -7, 1, -1, -6, 3, 10, 9, -13, 20, -13, -20, 7, -19, -62, -30, -17, -80, -48, -27, -12, -3, 42, 30, 37, 11, 33, 20, 78, 66, 40, 20, 14, -14, -15, 2, 20, 19, -1, -4, -40, 15, 53, -4, -4, -48, -70, -47, -31, 2, 48, 51, 13, -29, 39, 6, 9, -47, -13, -43, -26, -5, 41, -25, -9, -10, -18, -31, -70, -53, -20, -22, -60, -50, -38, -70, -81, -3, 2, 8, 52, 9, 18, 11, -5, -14, -29, -36, -40, -51, -45, -6, -8, -20, 10, -9, -2, -12, -13, -62, -47, -20, -48, -47, -33, -7, -15, -7, -3, -40, -19, -40, -7, -49, -42, -54, -48, -34, -34, -40, 4, 5, -16, -6, 37, 34, -4, -27, -18, -64, -48, -87, -57, -61, -81, -33, -18, -25, -46, -55, -37, -44, -36, -41, -89, -86, -76, -49, 15, -10, -1, -28, -22, 23, -29, -21, -24, -45, -53, -111, -73, -81, -61, -85, -60, -54, -63, -80, -44, -46, -14, -45, -56, -109, -161, -59, -7, 5, -14, -56, 6, 16, 1, -54, -25, -61, -57, -105, -81, -54, -49, -45, -31, -31, -29, -12, -33, -23, 0, -11, -20, -114, -129, -52, 16, -15, -46, -35, -48, 24, 5, -38, -31, -14, -40, -81, -44, -35, -1, 35, 42, 40, 24, 53, 34, 48, 23, 33, -12, -70, -91, 3, 11, 17, -65, 24, -99, 9, 41, -37, -14, -15, -26, -62, -43, 28, 47, 43, 57, 85, 79, 35, 51, 67, 51, 62, 34, -48, -98, 6, 5, -19, -83, -20, -66, 29, 13, -28, -41, -41, -24, 9, 24, 68, 69, 20, 10, 15, 38, 26, 81, 48, 58, 72, 15, -34, -41, -16, -42, -16, -55, -55, -54, -40, -4, -26, -31, -45, -19, 7, 51, 83, 71, 11, -15, 15, -14, 28, 59, 108, 86, 60, 16, 6, -29, -40, -29, 8, -57, -20, -9, -30, 25, 24, -38, -32, 16, 31, 66, 17, 35, 5, -22, -19, 1, 43, 28, 15, 43, 48, 33, 36, 35, 32, 23, 24, -31, -63, -33, -16, -7, 6, -26, -15, 10, 11, 67, 16, 34, -10, -15, -20, -4, 20, 16, 19, -4, 28, 108, 95, 44, 37, 44, 28, -41, -27, -18, 5, -8, -9, -16, 25, 22, 5, 5, 26, 36, -24, -31, 0, 10, -9, 43, 5, -13, 41, 96, 66, 31, 39, 47, 12, -61, 63, 15, -19, 53, 17, 33, 15, 24, -7, -19, 17, 44, -22, 4, 11, 36, 33, 30, 3, 22, 18, 33, 50, 25, 59, 62, 9, 20, 90, 41, 40, 29, 25, 32, 9, 27, 18, 21, 54, 45, 26, 18, 14, 22, 9, 23, 37, 48, 6, 26, 29, 8, 50, 36, 40, 16, 59, 51, 37, 12, 54, 45, 42, 63, 56, 41, 76, 75, 28, -1, 15, -15, -17, -19, 8, -11, -34, -10, 49, 16, 28, 47, 24, -2, 52, 25, 75, 44, 37, 36, 31, 53, 99, 62, 35, 5, 38, 0, -35, -59, -87, -19, -1, 1, 17, 26, 27, 35, 11, 72, 5, 6, 10, 58, 98, 91, 59, 63, 56, 32, 71, 38, 27, -4, -15, -43, -52, -53, -71, -24, 14, 62, 51, 75, 41, 33, 50, -1, -20, 1, 24, 108, 44, 104, 21, 27, -12, 5, -16, -2, 9, -8, -74, -63, -39, -34, -40, 8, 51, 50, 54, 69, 51, 35, 39, -46, -16, 12, 62, 59, 41, 9, 10, -6, -13, -22, -54, -17, -32, -35, -40, -55, 11, -26, 10, 38, 49, 20, 51, 57, 14, -23, 10, -16, -4, -18, -16, 38, 35, 23, 20, -25, -16, -46, -68, 3, -25, 9, 15, 11, 9, -2, -50, 23, 2, 42, 35, 32, -47, -17, -32, 12, 5, -34, 29, 69, 64, 50, -4, -2, -29, -30, -14, 8, 3, 28, 8, -9, -69, -66, -90, -56, -54, -34, -18, -42, -39, 28, -17, -17, 5, -13, 21, 35, 16, 0, 30, 1, -25, -49, -31, -14, -50, -39, -59, -122, -157, -140, -127, -170, -61, -72, -76, -64, 20, -18, 17, -8, 12, -20, -9, -49, -61, -115, -78, -100, -132, -213, -118, -102, -99, -91, -57, -63, -138, -159, -124, -128, -108, -80, -53, -42, -29, 7, 9, -11, -18, 2, -5, 6, -16, -39, -44, -52, -60, -64, -124, -130, -82, -22, -30, -74, -118, -92, -55, -68, -68, -68, -30, 6, -1, 16, 19, -16, 8, -6, 20, -18, 4, 3, 19, -15, 18, -6, -4, -20, 14, 15, -14, -1, 3, 4, 18, -13, -20, 20, -10, -11, 16, -17, -12, 20, 9, 907, 7, 12, 11, 19, -26, -5, -7, -5, -35, -18, -64, -16, 9, 17, -69, 8, -5, -52, -23, -1, -9, 16, -26, -6, 19, 0, -6, 2, -8, 1, -6, 30, 15, -44, -25, -53, -55, -15, 31, 51, 17, 6, -10, 58, 2, 5, 11, -1, 1, 32, 28, 88, -2, 5, 5, -13, -7, 4, 2, 12, 70, -11, 14, -15, -61, -38, 13, -13, -5, -3, 14, -5, 17, 54, 32, -34, -5, -24, -8, -51, -29, 19, 11, -7, -14, -8, -12, 28, 112, 50, 33, -11, 29, 34, -5, 32, 8, -9, -1, 25, 9, 28, 34, 11, -16, -52, -94, -29, -16, 3, -13, -9, 11, -26, 12, 56, 138, 79, 92, 73, 54, 19, -31, -3, -38, -46, 6, 21, 6, 43, 18, -4, -67, -72, -57, -11, 61, 8, -6, -19, 12, 11, 23, 32, 112, 128, 94, 41, 33, 22, -14, -15, -45, -27, -9, -8, 46, 2, -1, -1, -23, -8, -35, -5, 91, 26, 16, 5, 9, 43, 66, 98, 160, 120, 114, 59, 13, 39, 44, 9, 7, 1, 16, 10, 41, -20, 16, -23, -2, 15, 47, 33, 69, -19, -7, -7, -7, 20, 74, 72, 132, 139, 160, 113, 36, 67, 62, 40, 16, 24, 36, 26, 27, -11, 6, -32, -8, 46, 85, 41, 46, -15, -8, -8, -33, -14, 68, 83, 122, 148, 95, 54, 34, 60, 35, 28, 23, 20, 6, 29, 6, -4, -56, -19, 68, 92, 64, 15, 70, -55, -19, -7, 1, -11, 27, 115, 121, 96, 27, -3, 2, 13, 22, 5, 5, -1, -26, -4, -15, -14, 10, 44, 84, 124, 103, 83, 72, -57, -21, -20, 36, 34, 20, 33, 35, -9, -22, -50, -49, -37, -21, 28, 3, -26, -41, -33, -29, 23, 40, 90, 96, 93, 88, 91, 79, -13, -24, -17, -2, 6, 64, 48, 22, -39, -66, -51, -77, -56, -43, 7, 19, -28, -52, -5, 43, 104, 104, 54, 64, 87, 87, 58, 40, -31, -10, 0, 2, 0, 10, 37, -20, -52, -17, -70, -62, -33, 10, 37, 3, -44, -4, 49, 102, 129, 128, 74, 77, 69, 73, 13, 4, -44, 7, 13, -16, -72, -7, -16, -49, -2, -13, 18, -30, 14, 16, 20, 16, -6, 81, 169, 177, 121, 92, 41, 37, 14, -2, -13, -9, -97, -24, -11, -5, -48, -48, -22, 19, -3, 28, 0, 49, -3, 1, 36, -10, 32, 140, 236, 136, 68, 0, -33, 12, -15, -23, -66, -35, -84, -50, 11, -52, -47, -11, 28, 1, -1, 5, -31, 8, -14, -5, -11, -21, 8, 101, 114, 61, -34, -68, -77, -53, -26, -48, -69, -44, -60, -31, -23, -51, 20, 66, 140, 11, -39, -38, -40, 4, -14, 14, 32, -20, -15, -1, -4, -31, -119, -92, -41, -55, -33, -66, -45, -78, -66, -19, -32, -53, 25, 44, 63, 82, -30, -53, -62, 0, 19, 28, 2, -12, -25, -37, -26, -38, -81, -72, -40, -50, -71, -42, 6, -52, -39, -55, -48, -15, -2, 43, 27, 18, -27, -29, -13, -9, 2, 7, 15, 0, -26, -17, -3, 6, -45, -40, -35, -76, -69, -52, -28, -35, 2, -58, -46, -37, 5, 72, 55, -6, -54, -33, -19, -16, -16, -25, 32, 30, 4, 29, -8, 2, -16, -36, -64, -91, -52, -25, -44, -33, -3, -58, 34, 4, 3, 74, 17, -7, -26, -25, -39, -66, -48, -39, -8, 53, 38, 46, 54, 30, 44, 25, 27, -31, -17, -9, -43, -77, -27, -17, -7, -21, -22, 19, 44, 8, -18, -7, -3, -17, -18, 4, 8, 31, 42, 50, 50, 88, 81, 93, 65, 58, 4, -48, -57, -53, 24, 6, -3, 10, -6, -12, 26, 25, 53, 32, 67, 49, 33, 53, 17, 30, 9, 19, 43, 111, 102, 86, 68, 79, 45, 24, 25, 11, 11, -2, 16, -2, -21, 14, 12, -14, -17, -34, -4, -22, 31, 75, 35, 50, 79, 118, 124, 112, 135, 148, 95, 88, 120, 77, 21, -40, -42, -19, -7, 12, -14, -27, -11, -10, 24, 28, 15, -24, -15, -19, 33, 21, 70, 73, 95, 135, 129, 108, 126, 102, 55, 35, 8, 21, -19, 5, -1, 9, -5, 14, 6, 23, 26, 36, 27, 58, 10, 31, 23, 2, -21, 13, 62, 55, 87, 73, 25, 27, 23, 2, 29, 20, 2, 20, 18, -14, 6, -11, -20, 40, 24, 38, 32, -4, 20, 10, -17, -16, -3, 62, 45, 38, 40, 25, 24, 38, 32, -16, -9, 10, -12, -7, 7, 9, 20, 14, 10, -1, 1, -3, 5, -10, -11, -6, -5, 4, 3, -12, -1, 8, -13, -10, 17, 11, -8, 19, 15, -10, -17, 8, 18, -872, -16, 12, 18, 8, -9, 7, -11, 6, -34, -31, -11, 19, 23, 17, 12, -5, 15, 13, 18, 31, 32, 28, 10, -1, -18, -15, 0, 7, -3, 13, 4, 16, 5, 62, 32, 23, 20, 5, 29, 67, 71, 37, 70, 53, 68, 37, 18, -23, 0, 3, 24, 31, 6, 15, 5, -5, 9, -15, -36, 23, 54, 77, 49, 60, 28, 16, 49, 23, 30, 14, 58, 95, 48, 31, 72, 69, 30, 34, 45, 44, 30, 19, -10, -7, 13, -15, -58, -20, -11, 15, 6, 26, 11, -1, -36, -64, -15, -8, 13, -14, -13, -20, 14, -7, 20, 29, 36, 27, 47, -15, -4, 12, -19, 29, -15, 22, 7, 9, -13, -7, -50, -35, -40, -34, -20, -5, -24, -35, -22, 9, -24, -55, -49, 21, 23, 18, -7, -26, -13, -14, 3, 21, 10, 21, 43, 7, -18, 23, 3, -17, 3, -7, -18, 13, 0, 11, -12, 4, -15, -8, -38, -4, 17, 33, -25, -51, -21, 13, 9, -17, 5, 31, 24, 47, 27, 41, -11, 19, -6, 11, 12, 52, 6, 49, 20, 36, 23, 1, -12, -27, 30, 57, 15, -75, -33, 3, 0, -56, 17, 26, 49, 71, 47, 27, 27, 19, -5, -13, 19, 20, 20, 7, 13, 8, 53, 23, -23, -16, 17, 0, 27, -16, -19, 5, -28, -46, -20, 58, 52, 44, 35, 27, 13, -19, -9, 3, -9, 3, 10, 19, 47, -5, 9, 41, 19, 14, 18, 34, 47, 28, 30, -3, -54, -40, -37, -14, -8, 19, 19, 27, -12, -13, 14, 25, 5, -5, -19, -30, 1, -10, -20, 6, 7, 12, 18, 27, 71, -37, -14, -27, -89, -39, -83, -21, -15, 31, 42, 10, 10, 12, 15, -10, -10, -10, -13, -12, 3, 7, -31, 18, 27, 6, 6, -28, 28, -48, 22, 8, -32, -117, -94, -51, -56, 32, 18, 18, 5, 18, 5, 31, 0, 15, -15, 12, -11, -9, -36, 11, -19, -52, -43, -21, -34, -4, 24, 6, -30, -97, -104, -53, -54, -19, 38, 50, 31, 47, 39, 33, -1, -35, -19, 11, -27, 6, -5, 1, -3, -22, -9, -44, -69, -8, 27, 25, -37, -103, -93, -107, -92, -86, -5, 70, 46, 52, 18, 13, 2, -32, -23, -10, -26, 13, -18, -16, 13, 2, -52, -8, -26, 29, 6, 44, -42, -68, -96, -202, -166, -181, -133, -32, 23, 20, 22, 3, -4, -7, 9, 7, -12, -12, -24, -21, -15, 8, -32, -7, -23, -39, -5, 18, 11, -9, -90, -204, -277, -266, -295, -194, -73, -8, -18, -16, -38, -19, -37, -21, -24, -38, -12, -9, -22, -1, -44, -16, -30, -39, -16, -8, 28, 19, -45, -181, -274, -332, -329, -362, -262, -129, -97, -42, -45, -49, -46, -42, -51, -51, -6, -16, 1, -37, -13, 1, -16, -26, -29, 19, 22, 16, -20, -99, -181, -277, -284, -314, -367, -330, -241, -170, -102, -100, -24, -28, -18, -29, 6, 21, 15, -40, -47, -27, -27, -50, 0, -19, 24, 6, 7, -9, -69, -59, -65, -89, -128, -116, -143, -113, -53, -44, -36, -10, 3, -9, -18, 20, 26, -3, -54, -65, -62, -46, 1, 17, 8, 30, 53, 84, 77, 75, 77, 69, 33, 47, 20, 38, 24, 26, 5, 1, 42, -2, 8, 2, -5, -28, -10, -129, -30, -10, -1, -9, 26, 90, 120, 73, 74, 68, 92, 114, 99, 82, 70, 74, 57, 39, -4, 31, 2, 13, 2, -1, 1, -54, -49, -95, -71, -11, -18, -7, 2, 72, 135, 113, 37, 27, 37, 48, 75, 73, 65, 28, 48, 1, -26, 4, 5, 5, 2, -15, -26, -56, -66, -67, -49, -3, -5, 7, 24, 41, 69, 70, 78, 33, 11, 39, 7, 38, 47, 31, 14, 6, -2, -13, -9, -11, -4, -47, -111, -75, -15, -92, -15, -29, 20, -7, 26, 61, 70, 34, 74, 55, 54, 20, 3, 25, 25, 21, 4, -23, -27, -32, -35, -52, -58, -82, -51, -65, -50, -5, 23, -58, 3, 10, 18, 40, -10, -7, 16, 32, 73, 59, 40, 41, 18, 22, 52, 32, 0, -48, -54, -84, -54, -58, -36, -26, 5, 53, 31, 5, 20, 9, 12, -1, -25, -2, 39, 52, 21, 54, 64, 38, 68, 54, 47, 38, 45, 29, -14, -29, -54, -20, 59, 6, 14, 49, 18, 20, 7, 1, -19, -19, 0, 0, 10, 43, 56, 43, 52, 90, 61, 57, 52, 57, 84, 63, 43, 31, 48, 48, 42, 67, 26, 3, -20, -11, -8, 3, -16, -7, -15, 3, -13, -12, -12, 18, 12, 14, -17, -13, 4, -19, 6, 4, 12, -12, -14, 0, 14, -18, -9, 10, -17, -7, -3, 12, -1532, 4, 10, 18, -13, -4, -23, -6, 11, -40, -49, -3, -4, -24, -82, -69, -10, -18, -36, 4, 0, 4, -19, 1, -14, 16, 9, 1, 20, 14, -9, -3, -9, -26, 27, -17, -10, 28, -7, 29, 13, -7, -54, -44, -43, -58, -22, -84, -46, -80, -47, -66, -52, -15, 11, 10, 21, -1, 2, 26, 32, -5, -14, -25, -23, -23, -22, -27, -5, -31, -19, -2, 28, -30, 1, 5, 11, -15, -23, -41, -62, -12, 12, -11, -18, -7, 36, 41, 53, 4, 19, 6, -17, -42, 11, 12, -26, -51, -33, -18, -36, 11, 4, 20, 15, 31, 8, -1, 14, 24, -2, -11, 11, 8, 28, 30, 38, 39, 47, 20, 2, 4, -21, -25, -46, -25, -28, -13, 7, 4, 10, 29, 18, 25, 11, 48, 44, 62, 84, -15, -13, -17, 14, -3, 64, 83, 55, 66, 60, 45, 53, -7, -47, -22, -29, -41, -25, -9, -7, 2, -10, -4, 1, 2, 50, 37, 95, -12, 25, -6, 60, 41, 91, 91, 63, 78, 56, 71, 76, 38, 15, 5, -25, -24, -6, -14, 47, -3, 19, 36, 0, -1, 5, 87, 79, 37, 27, 17, 80, 95, 43, 53, 50, 56, 51, 20, 59, 42, 55, 17, 18, -7, 20, 37, 34, 25, 22, 17, 37, -33, -3, 43, 12, -9, -21, 36, 71, 124, 49, 12, 25, 53, 38, 32, 42, 63, 68, 54, 21, 33, 4, 26, 30, 43, 14, 9, 27, -9, -15, 66, -4, 1, -13, 35, 17, 92, 52, 4, -7, 13, 24, 10, 11, 23, 33, 17, 9, -45, -71, -40, -20, 1, -8, -18, -11, -8, -6, 77, -9, 30, 19, 26, 53, 66, 27, -3, -4, 9, -9, 24, 6, -5, -13, -18, 4, -52, -89, -79, -61, -89, -51, -28, 8, 15, 57, 96, 11, 38, -15, 70, 44, 53, 78, 28, 9, 21, 5, -3, -7, -19, -3, -46, -4, -25, -70, -59, -61, -62, -96, -28, -7, 59, 62, 89, 19, 44, 9, 49, 46, 44, 78, 8, -47, -14, -31, -11, -16, -17, 13, -28, -2, -21, -60, -24, 9, 2, -13, 32, 69, 46, 25, 57, -27, 1, 7, 39, 50, 30, -18, -17, -31, -21, -5, -34, -18, -21, -30, -1, 41, -2, 30, 17, 51, 84, 72, 65, 84, 22, -4, -4, -27, 0, 22, 1, 56, 6, -33, -82, -49, -25, -24, -30, -35, -8, -34, 4, 48, 67, 56, 68, 103, 72, 58, 17, -23, -65, -64, -34, -2, -12, -12, -21, 13, 20, -29, -51, -78, -45, -15, -43, 1, -14, 3, -23, 49, 42, 64, 65, 39, -39, -99, -140, -195, -119, -112, -52, -36, -32, 4, -30, 19, 31, 3, -59, -38, -56, -9, -33, -16, -5, -13, -27, -30, -44, -29, -62, -112, -214, -206, -210, -162, -107, -65, -65, -41, 11, 14, 11, 33, 62, -38, -21, -52, -34, -35, -18, -13, -17, -26, -62, -100, -122, -148, -165, -200, -200, -170, -166, -135, -83, -35, -13, 44, 23, 17, 52, 73, -14, -83, -61, 2, -50, -64, -49, -44, -14, -27, -65, -92, -113, -115, -145, -121, -74, -42, -58, -27, -6, 47, -24, 37, 0, -6, 4, 56, -48, -117, -61, -11, -53, -69, -49, -45, -20, -52, -16, -43, -21, -6, 10, 17, -9, 4, -2, 14, 14, 77, 9, -6, -1, -4, -21, 18, -45, -75, -42, 8, 8, 4, -8, 13, 23, -2, -7, 59, 31, 62, 79, 23, 52, 42, 35, 45, 26, 81, 29, -28, 74, -8, -28, 50, 28, -13, -10, -11, 11, 28, -7, 46, 27, 15, 4, 32, 57, 36, 58, 57, 15, -9, 27, 43, 20, 67, 53, -15, 17, -13, -11, -11, -8, 3, 17, 15, 4, 35, 0, 19, -6, 21, 11, -4, -2, 33, -3, 1, 1, 3, 19, 39, 76, 59, 70, 59, 14, 4, -32, -11, -6, 0, -36, -37, -41, -44, 2, 26, -7, 3, -6, -6, -21, 26, 3, 7, 23, 9, 20, 37, 64, 8, 31, 34, -15, 2, -14, -21, 19, -35, -92, -79, -43, -34, 21, 19, 17, -1, -7, -27, -3, 56, 16, 54, 43, 1, 23, 20, -1, 29, 16, 44, 18, -16, 18, 16, 31, 24, -12, -75, -74, -35, 14, 42, 9, 45, 32, 10, -10, 21, -21, 13, 6, -40, -61, -39, 0, -27, -12, 3, 20, 2, -20, 7, -5, -12, -17, -11, -52, -43, -69, -82, -27, 24, 21, 9, -43, -30, -37, -22, -28, -25, 14, -5, -9, -8, -15, 0, -14, -3, 3, -3, 12, 3, 13, 16, -4, -6, 5, 16, -10, -13, 13, -3, -15, -26, 9, -8, 5, -4, 13, -7, 17, 13, -14, 17, 0, -2, 110, -18, -13, -2, 14, 7, -3, -10, -32, 21, 10, 30, 2, 30, 55, 10, 1, -8, 21, -9, -3, 5, 19, 9, 15, 7, 4, 2, 5, -10, -10, 1, 8, 5, 6, 37, 27, 37, 35, 93, 58, -7, 4, -1, 54, 9, -14, -9, -24, -7, 1, 22, 39, 5, -5, 17, -8, -18, -8, 2, -7, 62, 71, 45, 16, 38, 42, 59, 43, 25, -8, -20, -11, 4, -14, -26, -9, -29, -55, -73, -65, 8, 2, -10, -4, -9, -22, -20, 17, 51, -6, -31, 21, 11, 51, 28, 25, -9, -4, 2, -26, -36, -3, -21, 8, -16, -26, -10, -55, -35, -49, 3, -17, -20, -24, -47, -57, 8, -11, -12, -5, -18, 24, 7, 20, -1, -8, -2, 4, -29, 10, -10, -4, -58, -7, 23, 27, -26, -71, -4, -14, -23, -22, -32, -5, 21, -25, -70, -1, 39, 26, 38, 14, 0, 8, -3, -4, 3, -23, -7, -34, -65, -44, -12, 1, -32, -127, -4, 13, -4, 12, -13, -24, -39, -59, -59, 15, -15, 43, 45, 2, -26, -32, -10, 8, 1, 15, 16, -53, -34, -5, 13, 6, -46, -96, -45, -4, 34, 12, -53, -15, -38, -69, -63, -16, 25, 38, 3, -32, -18, -45, -20, -19, 16, -7, -15, -4, -35, -12, 8, 8, -26, 14, 22, -11, -1, -20, -46, -59, -88, -89, -52, -6, 28, -7, 20, 2, -15, -20, -4, 42, 21, -24, -21, 1, -7, 20, 3, 12, -53, 20, 12, 3, 4, 10, -56, -121, -105, -104, -31, -17, 12, 20, 15, 14, 21, -2, -3, -2, -18, -41, -26, -4, 74, 52, 6, 42, -5, -53, -26, -34, 5, -39, -107, -79, -86, -60, -19, 16, 26, 33, 10, -5, 25, -3, -8, 7, 19, -23, -54, -9, 10, 48, 21, 12, 30, -74, -15, -19, -39, -114, -138, -107, -107, -99, -24, -1, 33, 16, -4, 2, -24, -21, -12, 30, 11, 1, -40, -11, -43, -5, 20, 33, 8, -56, 3, 0, -59, -112, -108, -136, -158, -122, -43, 0, -8, 47, 18, 11, -5, -11, -3, 36, 4, 21, 26, -16, -16, -46, -8, -40, -41, -35, -24, 4, -51, -97, -116, -124, -174, -178, -95, 41, -1, -1, -5, -7, -7, -27, 12, -10, 9, 29, 61, 5, -41, -62, -42, -53, -41, -27, 7, 34, -33, -104, -146, -201, -264, -276, -201, -58, 1, -40, -45, -25, -17, 19, 23, 31, 14, -5, 3, -26, 5, -57, -45, -66, -19, -16, 4, -4, -55, -50, -87, -176, -261, -345, -348, -248, -146, -74, -106, -104, -38, 17, 48, 39, 0, 17, 15, -42, -79, -91, -80, -71, -67, -4, -10, -22, -7, 35, -8, -15, -83, -195, -214, -270, -191, -128, -141, -90, -9, 7, 55, 9, -4, -3, -23, -83, -100, -108, -84, -59, -70, -24, -7, -1, -33, 34, 102, 109, 52, -29, -35, -83, -113, -107, -100, -24, 35, 36, 24, 42, 12, 31, -36, -85, -115, -132, -141, -107, -83, -60, 1, -29, -4, -7, 93, 130, 77, 58, 53, 19, -13, -34, -30, 2, 20, 26, 5, 17, 56, -10, -70, -98, -140, -115, -149, -91, -80, -63, -48, -2, -29, 8, 71, 118, 52, 50, 78, 56, 13, 4, -22, 14, 4, 4, 10, 24, 35, -19, -75, -98, -102, -112, -112, -89, -46, -53, -50, 5, 25, 52, 22, 0, 65, 35, 35, 48, 40, 6, -19, 2, 29, 61, 27, 34, 53, -21, -76, -131, -134, -154, -97, -98, -40, -34, -63, -7, 26, 43, 38, 52, 32, 32, 13, 56, 32, 22, -17, -3, 20, 40, 17, 34, 17, -51, -138, -170, -165, -128, -113, -63, -55, 14, -16, -9, 39, 27, 15, 29, 23, -36, -33, -14, 0, -17, -15, -30, -26, -2, -7, -18, -30, -89, -153, -153, -164, -116, -37, -73, -22, -17, 0, 19, 25, 3, 10, 27, 77, -12, -3, -17, -6, -1, -24, -35, -33, -30, -40, -64, -100, -174, -165, -162, -101, -97, -34, -18, -41, -21, 1, -12, 16, 62, -6, -1, 10, 40, 25, -2, -7, -12, -17, -48, -54, -58, -89, -89, -92, -115, -87, -80, -5, -6, -11, 51, 11, -28, -4, 1, -3, -15, 5, 2, 52, 95, 44, 38, 60, 58, 20, -6, -19, -9, 7, -45, -42, -57, -38, -46, -13, 8, 31, 57, 21, -4, -6, -20, 1, -2, -19, -6, 43, 62, 51, 38, 51, 52, 40, 41, 47, 38, 35, 51, -16, 1, -6, -22, 27, -4, 2, -7, -19, 13, -2, -19, 19, 8, 16, 10, -4, 7, -10, 14, 2, 7, -10, 1, 1, -4, -2, -13, -15, -4, -16, -13, -15, -2, -3, -10, -6, 6, -1, 12, -867, -14, -14, 13, 21, 30, 50, 41, 40, 12, 36, 51, 42, 80, 98, 33, 38, 39, 24, 38, 35, 56, 19, -2, 21, -10, -13, -17, 16, 17, 7, 17, -23, -37, 22, 57, 78, 42, 85, 97, 148, 171, 156, 104, 30, 53, 76, 87, 84, 101, 95, 32, 26, 3, 13, -11, -19, -2, -39, -33, 15, 46, 60, 87, 92, 76, 87, 53, 97, 63, 36, 25, 45, 7, 33, 65, 128, 84, 85, 91, 73, -12, 12, -9, 17, 17, -4, -41, -13, 66, 75, 74, 52, 10, 6, 85, 40, -9, -7, -40, -63, -37, -15, -20, 31, 74, 32, 54, 72, 81, 4, -20, -15, 1, -9, 13, 53, 53, 52, 59, 19, -12, 34, 14, -46, -40, -34, -62, -60, -47, -39, -49, -20, 25, -7, -45, -4, 14, -18, -3, -11, 7, -36, -22, 15, 37, 54, -2, 10, 2, 16, 27, -6, 15, -18, -60, -78, -58, -40, -33, -28, -34, -48, -42, -45, -1, 14, 21, 9, 16, -65, -28, 29, -9, 0, -19, -16, -2, 8, -3, 31, -8, -52, -43, -29, -46, -29, -61, -32, -18, -32, -38, -22, 37, 27, -13, -26, 13, -47, 25, 2, 23, 23, 8, 4, 14, 23, 31, 44, 4, -23, -25, -51, -40, -37, -3, -14, -26, -16, 26, 18, 59, -9, -34, 9, -32, -98, -44, -63, -33, -2, 12, 1, 28, 35, 46, 15, 8, -22, -42, -67, -45, -18, -27, -13, -5, -7, 34, 12, 24, -22, 6, 3, -2, 37, -93, -121, -16, 3, 14, -14, 22, 5, 63, 59, 22, -41, -44, -77, -16, -19, -30, -25, -5, -21, 16, -1, 50, 61, 18, 33, 23, -13, -91, -75, -13, 5, -4, 6, -7, 25, 60, 47, 12, -57, -50, -32, -29, -50, -51, -19, 11, -17, -1, 40, 9, 56, 24, 4, -20, -54, -213, -24, 13, 30, 6, 55, 12, 24, 43, 36, -11, -44, -58, -44, -68, -63, -67, -18, 13, 60, 75, 88, -1, 57, 39, 13, -25, -11, -137, -56, 10, 22, 25, 32, 30, 59, 87, 41, 49, -30, -43, -21, -31, -40, -14, -22, 54, 62, 83, 86, -20, 20, 26, -5, -22, -83, -84, -38, -20, 18, 27, 23, 44, 72, 82, 43, 27, -3, -29, 11, -27, 21, 17, 37, 51, 107, 58, 121, 11, 24, 38, -32, -51, -43, -30, -54, -47, -49, -32, -6, 12, 54, 50, 36, 0, -3, -14, -9, -4, 21, 27, 66, 39, 51, 43, 63, 5, 60, -17, 13, 9, -32, -90, -184, -51, -65, -41, -20, 29, 42, 34, 40, 6, 5, -36, -6, -6, 40, 24, 59, 11, 36, 47, 72, 36, 38, -3, 14, 37, -79, -30, -104, -74, -47, -20, 23, 29, 45, 47, 8, -8, -5, -6, -11, 2, 20, 7, 58, 14, 28, 48, 67, 60, 3, -11, -14, 40, -95, -13, -139, -32, 6, -4, 18, 25, 18, 48, 37, -13, -30, -26, -73, -51, -36, -19, 14, 52, 33, 22, 76, 53, 26, 8, 9, 25, -65, -84, -132, -77, -11, -7, 52, 57, 41, 37, 80, 56, 24, -17, -50, -82, -40, -37, -1, 16, 36, 90, 79, 55, 17, 37, 11, -26, -24, -141, -164, -112, -16, 13, 29, 56, 44, 76, 95, 85, 59, -20, -72, -67, -57, -46, -17, -1, 0, 79, 109, 71, 19, 0, -7, 3, -7, -84, -103, -81, -33, -2, 22, 64, 49, 84, 94, 60, 49, -17, -14, -51, -66, -7, 15, 18, 97, 134, 133, 102, 7, 36, 5, 19, -16, -52, -59, -101, -84, -21, 27, 23, 37, 35, 40, 22, -20, -12, -27, -14, 18, 52, 9, 55, 114, 116, 104, 73, 42, -13, -10, -15, -24, -62, -75, -106, -133, -138, -58, -13, 4, -14, -16, -16, -23, -15, -12, 9, 10, 29, 42, 77, 90, 137, 75, 23, -11, -18, 16, 3, 5, -53, -37, -159, -136, -122, -83, -32, 9, -39, -10, 5, 6, 22, 57, 49, 45, 10, 34, 67, 73, 64, 45, 31, 50, -12, 4, 12, -4, -33, -24, -110, -104, -71, 15, -39, -4, 42, 59, 66, 41, 27, 80, 107, 38, -23, 12, 10, 10, 26, -36, -27, -2, -10, -7, -8, 10, -6, -49, -68, -46, -91, -47, -27, -40, -15, -31, -64, -79, -91, -61, -72, -71, -115, -114, -56, -45, -20, -11, 18, -17, 13, -13, -11, 8, 9, -3, -36, -38, -52, -69, -65, -65, -79, -32, -54, -29, -37, -66, -45, -79, -35, -39, -15, -14, -15, -19, 2, 11, -11, -15, 7, 5, -17, -12, -11, 5, 13, -13, -15, 19, -11, 1, 12, 6, -1, -13, -4, 4, 16, 13, -10, -19, 5, 20, -13, 5, 3, 1, -1310, -5, 11, 15, 11, 20, 23, 36, 27, 39, 44, 69, -5, 1, -22, 41, -19, 1, 21, 5, 17, -16, 10, 11, 21, 16, -19, -19, 2, 14, 4, 11, -26, -32, 22, -16, -3, -19, 15, -39, -50, 3, -3, -28, -16, -50, -43, 18, -6, -2, -15, -8, -45, -27, -7, -3, 6, 14, -7, -2, -36, -4, -6, -50, -51, -73, -28, -58, -102, -49, -18, -39, -45, -40, -47, 22, 24, 29, -9, 71, 74, 27, -33, -16, 13, -6, 34, 31, -55, 2, 6, 15, -8, -15, -9, 3, -72, -67, -15, -30, -42, -10, -32, -13, 27, 27, 67, 87, -6, -44, -14, 17, 13, -13, 37, 16, -24, -27, -44, -83, -84, -26, -5, 44, 28, -4, -3, 8, 9, -45, -17, -2, -2, 57, 59, 42, -34, -74, -36, 15, 19, 9, 47, -33, -15, -37, -72, -69, -72, -24, -35, 19, 19, 14, 5, -60, -35, -68, 22, 22, 15, 26, -10, 25, -37, -94, -52, -20, 9, -19, 13, -46, -44, -69, -105, -90, -105, -100, -88, -72, -32, -16, -43, -61, -56, -41, -3, -4, -37, -21, -49, -27, -61, -138, -64, 10, -6, 9, 40, -49, -88, -117, -133, -101, -136, -166, -151, -112, -93, -49, -29, -42, -1, -1, -50, -80, -54, -59, -114, -104, -58, -110, -33, -14, -14, 41, 12, -47, -164, -170, -180, -148, -134, -169, -228, -155, -131, -108, -32, -10, -11, -1, -66, -77, -92, -76, -131, -126, -12, -4, 4, 35, 17, 42, 47, 6, -38, -85, -101, -38, -57, -96, -157, -163, -138, -72, 22, 17, 27, -37, -62, -75, -102, -137, -146, -102, -23, -53, 2, -5, 12, -55, 15, 19, -13, 8, 14, 31, 14, -9, -60, -82, -32, -2, 65, 58, 33, -4, -29, -37, -30, -80, -70, -75, -15, -71, -4, 20, -12, -54, -63, -60, -31, 30, 28, 88, 60, 6, -36, -1, 21, 47, 61, 43, 6, 1, -36, -26, 29, 11, -33, -52, -1, -11, -28, 15, 15, -1, 24, -16, -10, 89, 106, 79, 35, -16, -12, 23, 77, 66, 19, 34, 21, 9, -48, -23, 19, 5, -50, -25, 36, 20, 16, 22, -16, 3, -28, 6, 8, 73, 66, 55, 53, 4, -1, 10, 43, 62, 49, 24, 11, -11, -10, 0, 6, -13, -26, 34, 70, 89, 53, 5, -31, -37, 10, 10, -36, -30, 27, 54, -14, -41, -1, 0, 72, 76, 52, -2, 10, -5, -20, 10, 4, 9, 3, 20, 70, 97, 60, 35, 11, 43, 46, 1, -56, -89, -2, 11, -22, -21, -13, 23, 98, 123, 59, 20, 10, 0, -3, -31, 3, 13, -42, -30, 4, 80, 56, 58, 33, -3, -92, -83, -125, -82, -47, -10, -38, -2, -15, 19, 63, 108, 88, -12, 17, -20, 5, -40, 25, 30, 2, 25, -18, 42, 80, 53, 17, 6, -33, -51, -96, -88, -43, -13, -57, -27, -40, -17, 53, 116, 50, 28, -7, -22, -40, -16, -24, -10, 2, 19, 1, -26, 66, 47, 37, 2, -55, -71, -32, -44, -3, -17, -48, -40, 6, -13, 14, 69, 24, 20, 11, 5, -23, -3, -12, 24, 9, 14, 24, 7, 41, 70, -2, -31, -49, -28, -54, -1, 12, -14, -5, 1, 7, -11, -39, 21, 9, -6, 4, -17, -9, 20, 33, 6, 17, 7, 46, 43, 39, 49, -36, -7, 16, -53, -33, 19, -14, -18, 9, 7, 1, 26, -11, -56, -15, 4, -1, -18, -23, 20, -25, -2, 17, 4, 10, 49, 46, -21, -15, 10, 9, -90, -24, 2, 3, 16, -29, -35, 0, -17, -14, -12, -19, -5, 1, -7, -12, 3, -7, -2, -19, 10, -25, 10, 5, -14, -15, -45, -74, -75, -23, -34, -10, -54, -80, -104, -88, -88, -47, -10, -4, -52, 10, -2, -7, 33, 27, -28, -45, -2, -50, -5, 23, -10, 15, -66, -60, -100, -80, -16, -5, 13, -32, -16, -89, -101, -40, -63, -113, -59, -38, -22, -90, -100, -77, -69, -55, -26, -52, 0, 23, -6, 4, -12, -43, -67, -30, -38, -28, -51, -57, -66, -131, -92, -122, -159, -196, -174, -126, -137, -86, -86, -122, -83, -51, -19, -21, 2, 38, -18, -6, 4, 13, -24, -42, -45, -71, -87, -80, -70, -93, -88, -104, -109, -93, -79, -81, -60, -45, -22, -38, -54, -20, -26, -2, -16, -10, -8, -3, -1, -14, 4, 13, -26, -45, -27, -70, -24, -21, -58, -70, -45, 6, -53, -45, -61, -64, -23, -4, -21, -15, -9, -14, -10, 18, 12, 5, -19, 5, -2, 19, 2, -15, -4, -6, -2, 0, 0, 8, -1, -9, 1, -23, 4, 17, -6, -7, 7, 11, 1, 0, 16, 15, -13, 9, -1619, -7, -12, 5, -19, 1, -23, -36, -12, -25, 36, 39, 14, -16, -12, 60, 9, -6, 39, -5, 33, 15, -16, 30, 35, 15, -20, -10, -21, 3, 7, 9, -21, -41, -41, -56, 10, 25, -7, -16, -5, 8, -28, -3, -57, -27, 17, -15, -28, -48, -64, -15, -103, -31, -18, -16, 19, -12, 3, 11, 49, -41, -40, -64, -60, -3, -35, -44, -42, -21, -20, 9, 24, 23, 5, 22, 41, 5, -17, -17, 8, 7, -2, 4, 10, 7, 20, 23, 29, -31, -58, -69, -114, -77, -56, -28, -30, -9, 35, 10, 8, 11, 17, 32, 64, 29, 22, 22, 6, 56, 15, 20, 16, -13, 28, 2, -10, -8, -42, -61, -49, -62, -34, 13, 22, 0, -19, -5, 18, 65, 66, 67, 28, 63, 75, 9, 18, 7, 31, 21, -12, -4, 38, -2, 27, 0, 19, -14, -10, -6, 12, 5, -3, 29, 19, -13, 12, 31, 27, 16, 48, 33, 56, 15, -44, -17, 75, -17, -13, -17, 45, 73, 62, 33, 1, -10, -17, 11, 27, 14, 31, 35, 22, 17, 22, 3, 10, -2, 42, 36, 40, 21, 17, 3, 49, -8, -19, -10, 52, 34, 24, 21, 25, 9, 12, 10, 42, 54, 57, 7, 17, 12, 1, 25, 11, 13, 58, 55, 61, 50, 75, 56, -18, 1, 9, 32, 36, 71, -5, 17, 23, 36, -6, -10, 5, 51, 39, 42, 31, -17, -30, -23, 32, 34, 27, 42, 38, 42, 67, 75, 22, 48, 8, 16, 81, 80, 37, 5, 25, 9, -17, -15, 12, 34, 24, 35, 1, -46, -23, 9, -25, -26, -4, -5, -31, 32, 70, 27, -4, -2, 34, 24, 90, 67, 53, 39, 19, 15, -31, -13, 0, -8, -11, 22, 5, -27, -2, -41, -17, -18, -7, -51, -32, 34, 18, 41, -6, 29, 4, 32, 75, -1, 42, 20, 28, 26, -14, -9, -15, 0, -2, -10, 10, -1, 10, -17, -24, -22, -28, -25, -43, -45, -2, 21, 3, 27, 21, 19, 38, -21, 8, 10, 13, 13, -3, -48, -16, -11, -26, -13, -15, 2, -45, -60, -33, 3, -47, -52, -25, -17, -14, -14, 46, 3, -2, -18, 68, -4, -25, -66, -92, -34, -57, -21, 3, -28, -7, -21, -18, -31, -56, -80, -44, -58, -64, -47, -70, -87, -47, -40, 22, -20, -20, 17, 51, 1, -85, -152, -146, -111, -51, -40, 5, 25, -44, -61, -8, -40, -76, -81, -74, -82, -59, -87, -83, -95, -75, -34, 21, -18, -10, 5, 77, -4, -123, -189, -126, -71, -28, -46, -17, -37, -15, -39, 2, -35, -62, -93, -70, -95, -64, -72, -58, -62, -58, -57, -1, 1, 19, 0, 39, -8, -110, -101, -56, -41, 0, 12, -10, -9, 14, 9, 24, 1, -80, -97, -91, -114, -69, -43, -32, -32, -27, 25, 17, 64, 29, 24, 44, 68, -82, -61, -25, 13, 51, 38, 24, 65, 60, 88, 118, 101, -16, -81, -71, -65, -54, -19, -10, 6, -1, 15, 54, 45, 31, 49, 11, -19, -61, 4, 56, 38, 49, 48, 54, 34, 69, 91, 140, 104, 19, -40, -43, -38, -19, 21, 29, 5, 37, 19, 45, 51, 16, 7, 3, -41, -84, 7, 64, 39, 40, 53, 45, 37, 24, 39, 75, 78, 30, 4, 3, 4, 23, -11, -20, 11, 61, 19, 1, 26, 14, -3, 3, -94, -64, 26, 33, 29, 27, 6, 18, -13, 13, -15, 41, 45, 43, -4, -20, -36, -10, -24, 10, 13, 84, 98, 18, 68, -18, -7, -16, -110, -56, -3, 3, 20, -7, -7, 4, -9, 27, -7, 51, 47, -3, -6, -14, -25, -23, -24, 21, 41, 36, 75, 8, 32, 12, -23, -36, -81, -90, -30, -16, -11, -1, -3, -6, -5, 30, 37, 53, 52, 8, -23, -17, 7, 23, 42, 31, 43, -7, 42, 7, -9, 9, -30, -51, -57, -81, -78, -60, -46, -29, -1, 8, -10, 7, 48, 35, 53, 20, 35, 29, 8, 9, 22, 23, 2, -15, 57, 13, 1, -14, 17, 1, -24, -67, -110, -92, -49, 6, 7, 22, 34, 65, 34, 14, 24, 43, -3, -2, -17, 11, 6, -13, 9, -3, 11, 16, -17, 11, -3, 18, 35, 6, -28, -51, -11, -28, -20, 32, 16, 25, -34, -27, 15, 17, -12, 5, 11, -17, -52, -30, -21, -20, 25, 20, -14, 6, 20, 5, -14, 2, 0, -3, -23, -67, -37, -41, 12, 28, -20, 7, 18, -1, 12, -44, 2, -10, -9, -36, -8, 17, -12, 18, 5, -6, 21, -13, -6, -12, -6, 18, -19, -4, -15, -7, 17, 8, 15, 26, -9, -2, 12, -11, -15, -10, -7, 5, -16, -2, -8, 10, -19, 3, 1112, -16, -3, -19, -19, 5, 55, 36, 15, 33, 65, 42, 35, 50, 99, 76, 50, 55, 55, 46, 23, 18, 6, -12, 23, -6, -9, -14, 6, 8, -7, -7, 9, 25, 15, 58, 33, 69, 83, 88, 48, 108, 137, 154, 156, 84, 122, 102, 81, 140, 89, 75, 62, 9, -9, 1, 13, -7, -19, -2, -12, 5, 22, 78, 57, 85, 81, 174, 200, 172, 149, 151, 157, 189, 168, 97, 102, 125, 96, 100, 82, 25, -8, -13, 16, 4, -37, -67, -27, 12, 31, -4, 69, 45, 52, 51, 155, 103, 78, 63, 30, 60, -6, -1, 29, 63, 52, 24, 76, -3, -9, -1, -3, 17, -57, -50, -59, 9, 53, 10, 11, 48, 82, 51, 83, 51, 37, 58, 45, 23, 0, -7, 0, 5, 19, -22, -18, -2, -78, -4, -10, -4, -42, -44, -8, 10, 31, 27, 0, 1, 31, 26, 45, 2, 37, 9, 43, 37, -37, -50, -17, 12, -1, -36, -39, -54, -35, 3, 11, 6, -39, -78, -58, -4, -9, 6, 3, 6, -31, -42, -37, -31, -22, -3, -13, 4, -53, -35, -25, 2, -9, -28, -51, -135, -39, -14, 3, 1, -37, -22, -48, -27, -22, 12, -2, -2, -55, -47, -101, -80, -80, -28, -39, -42, -45, -32, -53, -7, -42, -25, -82, -131, -57, 14, -7, -50, -10, -108, -60, -37, -26, -26, 20, 27, -39, -86, -94, -109, -100, -71, -48, -47, -41, -37, -25, -24, -39, -66, -69, -110, -37, -28, -16, -31, 41, -115, -47, -42, -60, -30, 45, 23, -55, -53, -89, -76, -59, -51, -45, -11, -21, -13, -29, -8, -18, -24, -71, -106, 4, 10, 44, -29, -16, -82, -18, -39, -62, -47, -17, -44, -59, -34, -67, -19, 2, 18, 11, 6, 14, 23, 37, 13, -25, -64, -98, -85, -26, -36, -1, -68, -63, -101, -67, -50, -78, -83, -20, -49, -35, -35, -26, 18, 19, 26, 33, 1, 58, 58, 68, 9, -15, -88, -76, -70, -51, -27, -11, -39, 8, -46, -96, -73, -22, -26, -14, -31, 3, 13, -7, 30, 27, 22, -3, 26, 21, -3, -4, 1, -49, -56, -28, -28, -32, -31, -23, 27, -12, -30, -77, -51, -65, -25, 18, 34, 11, 27, -2, 40, 22, -3, -29, -9, -53, -80, -25, -26, -47, -41, 38, -29, 38, 42, -4, -19, -9, -3, -44, -32, 7, 17, 49, 10, 6, -2, 14, 44, 22, -3, -50, -35, -73, -37, 15, 8, -24, -5, 68, 36, 51, 38, -26, -1, 41, 24, -1, 1, -14, 32, 27, -11, 3, 2, 29, 15, -30, -3, -51, -29, 20, 53, 24, 28, 35, 34, 29, 83, 100, 34, -10, 21, 79, 19, 28, -10, 3, 13, -7, -53, -23, 6, -12, -15, -15, -6, -17, 19, 70, 81, 79, 38, 37, 50, 51, 7, 49, -47, 0, 50, 1, -1, -9, 2, -8, -2, 26, 35, 11, -13, -36, -59, -42, -29, 26, 43, 68, 74, 31, 6, 30, 0, -12, 1, 44, -4, -5, 3, 24, 32, 32, 49, 41, 39, 3, 59, 51, 13, -29, -51, -41, -27, 41, 88, 93, 105, 17, 14, 70, 31, -46, 1, 84, 27, 21, 39, 14, 42, 83, 60, 63, 55, 18, 61, 43, 7, 32, -38, -38, 5, 39, 70, 75, 96, 59, 89, 70, 44, -7, 12, 59, -20, -21, -33, -21, 7, 38, 48, 57, 53, 47, 26, 26, 57, 49, 24, -28, 2, 40, 42, 80, 66, 90, 69, 48, 37, -32, 22, 20, -4, -3, -12, -32, 5, -11, 33, 31, 32, 43, 23, 33, 57, 45, 32, 3, 13, 35, 21, 69, 63, 85, 46, 35, -6, -71, -35, -15, -10, 20, -24, -30, 63, 5, -13, 20, 20, 4, 19, 24, 51, -7, -21, 6, 2, 75, 44, 6, -6, 14, 7, -17, 14, -57, -36, -26, -3, -18, -21, 62, 86, 108, 46, 23, 9, -6, 27, 39, 48, 5, 4, 10, -13, 11, -28, -62, -79, -81, -49, -71, -36, -43, 13, -8, -13, -5, 5, -31, 2, 38, 47, 90, 60, 15, 31, 63, 31, -9, -69, -78, -121, -140, -121, -143, -169, -167, -89, -67, -41, -51, -61, -8, 13, -2, 16, -18, -13, -32, -58, -45, -26, -49, -55, -6, -38, -46, -84, -62, -108, -137, -132, -67, -83, -46, -54, -18, -34, -10, -37, -1, -17, 14, -16, -20, 15, -4, -43, -30, -41, -55, -45, -39, -14, -42, -47, 17, -1, -48, -61, -55, -33, -24, -21, -37, -3, -22, -16, -11, -19, 13, 5, -5, -12, 6, -15, 4, -14, 8, 6, 16, 14, -15, -11, -10, -25, -19, -20, 10, 15, -10, -1, 0, -13, -19, -14, 15, -2, -3, 76, 2, -16, -19, 11, 36, -31, -47, -41, -46, -48, -70, -85, -100, -122, -24, -20, 1, -34, -14, -39, -25, -18, 25, 17, -13, -17, 7, -11, 20, 8, 22, -8, -17, -73, -86, -90, -113, -145, -136, -130, -111, -215, -139, -116, -174, -154, -159, -119, -90, -58, -34, 5, 4, 14, 19, 16, 8, 5, 6, -8, 17, 11, -41, -46, -88, -67, -58, -50, -44, -40, -71, -58, -67, -79, -36, -89, -53, -61, -17, 17, 24, -9, 18, -15, -6, 49, 36, -35, -52, -7, -2, -17, -13, -32, -18, -39, -35, -1, -23, -75, -36, -12, -7, -13, -46, -47, -30, -52, -41, -23, -3, -2, -3, 81, -10, -63, -77, -37, 22, -28, 0, -22, -44, -68, -58, -48, -75, -37, -45, -14, -40, -81, -66, -52, -18, -21, -42, -3, 14, -10, -18, 36, -6, -54, -73, -11, 23, -9, -5, -28, -65, -55, -74, -109, -82, -98, -86, -16, -51, -83, -134, -128, -42, -21, -6, -7, 1, 28, 6, 50, -26, -11, -44, -21, -31, -69, -48, -20, -36, -35, -52, -59, -57, -62, -72, -26, -31, -61, -100, -89, -67, -27, -21, -27, 9, 16, -12, 34, -14, -38, -38, -45, -35, -43, -54, 4, 35, 4, -2, 33, -19, 17, 17, -5, -13, -9, -9, -14, -54, -7, 2, 13, -27, -10, 20, 20, 29, -28, 14, -58, -29, -29, -14, 36, 9, 48, 49, 78, 80, 35, 24, 28, 37, -6, 9, 27, 25, 45, 47, -16, -15, -14, 34, -21, 64, 74, 26, -13, 36, -26, -3, 29, 27, 44, 64, 58, 61, 69, 28, 10, 36, 7, 12, 16, 54, 49, 36, -3, 19, -40, -12, -14, 59, 30, 40, 37, 65, -8, 12, 53, 16, 40, 38, 68, 80, 21, 12, 27, 27, 48, 40, 90, 93, 30, -21, 7, 12, -2, 26, 47, 66, 64, 0, 42, 33, 23, 10, 33, 27, 53, 56, 63, 63, 40, 30, 29, 45, 67, 36, 92, 82, 41, 40, -2, 17, -24, 23, 41, 18, 15, 25, 34, 25, -38, 20, 18, 35, 15, 44, 39, 67, 46, 39, 22, 29, 65, 49, 62, 78, 76, 54, 20, -5, 24, -4, -9, 55, 35, 46, 76, 11, -6, 13, 11, 29, 48, 28, 25, 27, 66, 26, 50, 35, 64, 41, 51, 97, 56, -12, 6, -22, 21, -7, -21, 25, 61, 52, 89, 76, 24, 5, 35, 10, -10, 25, 37, 47, 73, 85, 45, 45, 29, 8, 28, 40, -7, -50, 3, -20, 23, 6, -15, -20, 18, 16, 39, 31, 1, 7, 13, -43, -17, 2, 41, 108, 129, 83, 54, 40, 33, 9, -13, -20, -13, -26, -15, -1, 8, -17, -39, -1, -29, -5, 38, 33, 15, 38, -6, -18, 40, 52, 108, 92, 105, 37, 14, -7, 2, -15, -23, 3, -27, -65, -30, -1, 1, -2, -16, 41, 11, 41, 50, 41, 28, 22, -17, 28, 55, 118, 115, 90, 64, 11, -26, -40, -58, -33, -85, -4, 14, -58, -40, -9, -14, 27, -71, 2, 31, 42, 53, 29, 21, 14, 27, 34, 88, 90, 28, 18, -18, -58, -80, -56, -55, -80, -61, 10, -12, -58, -3, -18, -30, -42, -51, 40, 51, 28, 44, 21, 8, -15, 4, 34, -20, -28, -87, -89, -117, -63, -43, -50, -90, -65, 1, 1, -6, -32, 6, -4, -2, -17, 9, 32, 46, 26, 9, -27, 12, -12, -25, -34, -102, -158, -145, -119, -102, -73, -82, -66, -82, -42, -12, 28, -3, -37, -29, -34, 14, -16, -12, -40, 6, 30, -28, -32, -66, -67, -94, -135, -119, -161, -155, -120, -91, -66, -66, -84, -103, -85, -12, 32, -11, -63, -26, 12, 3, 1, -37, -52, 0, 36, -29, -37, -45, -91, -109, -86, -92, -35, -52, -88, -42, -76, -14, -28, -12, -29, 32, 56, 9, -43, 44, -1, 16, -15, -53, -39, 8, -8, -16, -24, -38, -27, -81, -83, -96, -68, -31, 31, 15, -23, -8, 0, 2, 12, -6, 28, -25, -56, 17, -13, -11, 18, -32, -42, -45, -40, 23, 17, -43, -8, -74, -65, -78, -36, -42, -36, -47, -29, 3, 43, -5, -30, 6, 15, 1, -26, 6, -4, 7, 3, 7, -2, 6, -6, -40, -9, -27, -17, -45, 23, -11, 26, 34, 25, -5, -9, 32, 64, 18, 24, 35, -2, 4, -22, -10, -10, 12, 17, -13, 7, 11, -30, -17, 2, -43, -36, -56, -46, -49, 5, 1, -49, -21, -16, 3, -20, -9, -32, -9, -3, 19, -12, 20, 2, 18, -18, 19, 17, -2, 18, -17, -15, 20, -4, -5, 15, -9, 18, 16, 7, -12, -17, -7, 5, 15, -6, 14, -10, 12, 20, 4, -3, 5, 1160, -15, 12, -2, -2, 22, 43, 4, -24, -16, 8, 33, -26, -49, -66, 20, 2, -26, -4, -17, -15, 5, -5, 17, 0, 0, 3, 3, 1, -5, -20, -11, -12, 33, 35, 15, 3, 40, 5, -19, -25, 10, -76, -18, -14, -11, -34, -60, -51, -71, -101, -50, -55, -16, -17, -16, 13, -11, -4, -5, 26, 27, 54, 45, 13, 63, 15, 36, -2, -3, -13, 20, 56, 39, 15, 57, 5, 5, -15, 23, 43, 17, 4, -12, -17, 4, 38, -10, 26, -26, 2, 29, 22, 1, 24, 39, 0, 20, 20, 26, 37, 39, 45, 81, 30, 43, 39, 64, 94, 93, -4, -14, 18, 6, 17, -25, -9, -27, -11, 31, 42, 10, 27, 35, 18, 16, 12, -25, 10, 43, 54, 54, 10, 4, 13, 90, 104, 78, 37, -18, 3, -8, 13, -47, -26, 3, 21, 37, 22, 24, 11, 25, -18, -1, -13, -10, 5, 28, 0, -8, 21, 25, 35, 48, 30, 18, 9, 15, -7, 14, -27, -40, -2, 18, 24, 47, 41, 34, -3, -25, -44, -19, 9, 6, 26, 35, -11, -20, 13, 12, 18, 50, 21, 15, -12, 5, -16, -2, -17, -89, -30, 46, 30, 24, 28, 19, -8, -5, -28, -19, -31, -35, -11, 2, -39, -5, 9, -10, 13, 29, 7, 6, 35, 23, 3, 5, -52, -43, -17, 25, 48, 31, 24, -34, 10, -9, 13, -27, -30, -2, -45, -83, -80, -68, -53, -8, 25, 33, 47, 27, 26, 62, -16, -19, -40, -66, 0, 21, 37, 37, 30, -9, -8, -4, 2, -23, -62, -68, -89, -90, -110, -137, -69, -28, -24, -10, 13, 15, 16, 30, 22, 2, -34, -69, 32, 58, 3, 9, 17, -9, -10, 17, 8, -21, -92, -104, -49, -38, -31, -65, -66, -68, -49, 14, -17, 22, 1, 26, -18, 25, 21, -4, 85, 45, 1, -12, -20, 2, -14, -14, -22, -33, -53, -59, -25, -32, 26, 9, 12, -18, -39, -9, -48, 8, 39, 22, -12, 13, 19, 6, 94, 49, -18, -3, -54, -50, -25, -35, -29, -25, -38, -42, 3, -17, 46, 65, 58, 63, 16, 6, -14, -18, 53, 25, 30, -2, -29, -7, 76, 31, -46, -48, -77, -130, -93, -54, -50, -20, -26, -12, -22, 12, 44, 63, 56, 70, 27, 16, -10, -4, 51, 7, 5, -37, -16, -7, -17, -72, -112, -106, -103, -125, -66, -63, -76, -73, -10, 25, 41, 37, 48, 60, 27, 13, -6, 32, -37, -29, 36, 9, 5, -40, 57, 30, -64, -101, -109, -142, -136, -98, -92, -85, -117, -104, -27, 27, 49, 51, 59, 1, -13, -9, 9, -4, -20, 13, 32, 12, -16, -14, 77, 113, 23, -10, -36, -51, -50, -22, -25, -51, -79, -66, -34, 11, 33, 27, 34, -6, -52, -73, -17, 10, 1, 26, 75, 19, -1, 4, 107, 138, 128, 76, 19, 45, 31, 31, 55, -3, -29, -25, 7, 59, 46, -5, -12, -32, -39, -58, -1, -28, -4, 30, 66, 6, 42, 46, 22, 161, 140, 72, 43, 58, 31, 72, 91, 65, 47, 22, 35, 30, 9, 5, -24, -12, -26, -10, -10, -9, -9, -61, -18, 13, 39, 1, 37, 57, 108, 75, 33, 44, 53, 64, 57, 28, 36, 21, 8, 25, 21, -7, -10, 11, -2, -23, -4, 25, -62, -45, -18, 29, 10, 62, 49, 32, 8, 41, 28, 36, 7, -6, 17, -6, -12, -21, 4, 7, -13, 29, 6, 20, -26, 10, 24, 12, -13, -35, -2, 54, -3, 34, 54, 14, 52, 18, 2, 18, 8, -10, -17, -16, -40, -4, -1, 16, -1, -23, 3, -44, -28, -22, -7, 38, 27, -6, 35, 26, -9, -6, 56, 31, 26, 49, 1, -20, -41, -56, -95, -63, -31, -69, -23, -24, -32, -43, -35, -37, -1, -26, -28, -10, 4, -10, -9, 8, -13, -46, 39, 37, -13, -34, -18, -36, -75, -87, -53, -66, -45, -22, -46, -36, -31, -13, -37, -39, -58, -34, -74, -27, -19, 20, -12, 12, -8, 18, 41, -13, -63, -75, -42, -34, -12, -49, -5, -18, -56, -33, -39, -66, -32, -40, -81, -93, -4, -35, -10, -22, 11, 3, -18, -13, 1, 21, -13, -15, 5, -1, 0, -8, -18, -2, 21, -7, -34, -84, -107, -91, -67, -51, -81, -29, -13, -7, -21, -23, 20, 15, -9, -19, -14, -10, 0, 18, 2, -12, -12, 14, -22, -9, -10, 0, 5, -47, -28, 3, 12, 15, -2, -21, -17, -23, 15, 12, -15, -14, -16, -10, -9, 4, 21, -1, -17, 12, -8, 3, -2, 19, 20, -1, 2, -18, -6, -1, -2, 6, 14, -11, 12, -15, 1, -3, 4, -3, -10, 19, -19, 1827, -13, -3, -14, 1, -30, -29, -6, -18, 0, 3, -40, -46, 7, -24, -85, -13, -4, -51, -50, -19, -14, -9, -35, -6, 10, 15, 9, -9, 2, -15, -3, 5, 29, -39, 35, 2, -43, -8, -16, -74, -62, -39, -7, 24, 17, 5, 28, -5, 1, 41, 41, 75, 21, 7, -9, 14, -13, -13, -31, 14, 70, 20, 16, 30, 61, 16, 4, 0, -21, 19, 19, -6, 25, 63, 28, 5, 49, 11, -2, -58, -28, 61, 5, 20, 8, -8, -47, -43, 69, 8, -22, 39, 42, 25, -16, 40, 7, 31, 59, 43, 64, 71, 55, 83, 60, 35, -18, 52, 70, 24, -17, 10, -10, 10, 9, 22, 61, 33, -25, -11, 26, 4, 11, 39, 24, 0, 11, -3, 1, 1, 44, 62, 57, 28, 14, 64, 109, 38, -16, 12, 11, 34, 14, -22, -17, -49, -45, -32, -39, 8, -2, 4, 19, 6, -18, 4, 2, -19, -29, -32, 4, 3, -27, 81, 54, 12, 23, 1, 12, -37, -18, -45, -75, -23, -58, -47, -31, -9, 25, 16, 26, 13, -17, -40, -66, -65, -79, -38, -21, -14, -27, 41, 36, 40, 33, -4, 23, -61, 36, -25, -50, -4, -27, -20, -27, 14, -9, 5, 14, 14, -25, -64, -100, -86, -101, -91, -72, -60, -60, -39, -4, 19, 18, 12, -14, -55, -20, 15, -25, -45, 0, -47, -30, 9, -2, -5, 12, -27, -24, -41, -78, -85, -75, -100, -98, -99, -88, -89, -16, 6, -1, -10, -51, -58, -52, -1, 7, 4, -27, 0, -51, -60, -33, -25, -6, 42, 47, 38, 2, -33, -63, -53, -82, -65, -77, -99, -66, 9, 21, -22, -40, -44, -42, -1, 25, 37, -2, -26, -18, -35, 13, -12, 38, 65, 71, 70, 81, 37, 36, -11, -32, -66, -140, -110, -32, 1, 36, 3, -47, -38, 16, 25, 64, 47, -50, -44, -21, -3, 30, 21, 15, 89, 83, 105, 100, 58, 68, 26, -20, -19, -86, -131, -28, -14, 9, -25, -61, -19, 30, 43, 56, 86, 0, -15, 34, 41, 53, 45, 2, 51, 85, 93, 83, 96, 61, 54, -24, -51, -68, -51, -21, -27, 42, 12, -35, -11, 40, 59, 98, 64, 20, 18, 50, 37, 49, 28, 45, 39, 74, 98, 96, 68, 64, 6, -25, 0, 5, 24, 1, -16, 36, 10, -6, -14, 27, 69, 115, 67, 50, 32, 45, 43, 41, 32, 53, 97, 103, 113, 97, 54, 5, 18, -23, 29, 72, 122, 67, -14, 31, -17, 5, 28, 17, 55, 100, 40, 27, 6, 32, -11, 2, -4, 72, 160, 202, 110, 58, 19, -9, -35, 8, 31, 81, 88, 40, -1, -26, -35, 17, 46, 29, 65, 49, 15, -39, -18, -7, -13, -34, -14, 57, 166, 170, 105, 21, 3, -20, 16, 41, 37, 63, 86, 40, -15, -55, -28, 27, 37, 41, 43, 19, -43, -53, -38, -32, -53, -111, -100, -3, 95, 79, 69, -6, -30, -42, 5, 45, 21, 6, 50, 20, -36, -55, -23, 28, 119, 108, 0, -18, -54, -41, -39, -69, -104, -124, -127, -43, 48, 41, 28, 0, -12, -22, 9, 19, 6, 6, 16, 26, -6, -73, -43, 14, 95, 98, 56, -38, -69, -19, -53, -53, -70, -84, -69, -59, -21, 35, -19, -7, -33, -9, -1, 19, 24, 33, 23, 13, 10, -69, -4, 4, 67, 71, 15, -76, -72, -72, -65, -74, -46, -49, -48, -7, 2, 6, -20, 3, 0, 3, 11, 8, 7, 47, 44, -42, -9, -47, -13, 33, 80, 105, 12, 0, -51, -54, -21, -51, -50, -38, -3, 19, 23, 9, 11, 9, -7, 20, 2, 21, 19, 21, 55, 25, 11, -6, -13, 56, 84, 68, 15, -18, -25, -36, 18, -9, -10, -27, -15, -4, 5, -13, 25, 4, -16, -23, -37, 5, -2, -13, 51, -13, 25, -1, -8, 30, 69, 62, 80, 82, 23, 27, -16, 2, -56, -52, -33, -16, -6, -6, -27, 6, 4, -3, 7, 2, 16, 34, 56, 5, -48, -14, 6, 1, 26, 63, 84, 123, 55, 54, 37, 6, 9, -12, -65, -35, -18, -47, 4, 38, 59, 62, 65, 50, 33, 43, 32, 5, -28, -10, -5, 17, -13, -28, 26, 42, 32, 24, 26, 17, 11, 7, 5, 12, 16, 28, -1, 42, 58, 24, 12, 13, 27, -7, -10, -21, 0, -15, 5, 19, -6, 11, -4, -4, 12, 54, 51, 49, 45, -2, -12, 22, 39, 18, 28, -9, 37, 22, 45, 29, 28, 1, 7, 5, 16, -13, 0, -16, 1, -11, 18, -19, 0, -8, -7, 8, -4, 4, 4, -7, -3, -9, 18, -16, 7, -18, 15, -16, 1, -8, 5, -6, 20, -12, -20, -2546, 14, 18, 1, 12, 1, 11, 17, 5, -19, -38, -7, -9, -44, -74, -48, -33, -32, -3, -19, -14, -7, -3, -17, 7, 12, -18, -8, 3, -9, 10, -14, 3, 7, -18, -23, -4, -23, -6, 21, -10, -39, -87, -62, -52, -54, -44, -60, -46, -88, -70, -67, -44, -10, -6, 15, -1, -5, 24, 2, -12, -74, -53, -25, 15, 47, 29, -2, -25, -31, -13, 17, 13, -54, 14, 30, 23, 2, 27, -13, 0, -22, 18, -15, 19, 12, 34, 28, 58, -38, -10, 44, 14, -13, -2, 15, 14, -16, 7, 10, -21, -22, -9, 4, 18, 2, -30, 13, 36, 51, 33, 2, 13, -18, 15, -35, 8, -24, -44, 10, -4, 1, 4, -14, -17, 14, -35, 1, -23, -22, -3, 16, 5, 15, -11, 16, 43, 75, 47, -11, 13, 7, -27, -20, 23, -66, 8, -13, 13, 21, 9, -24, -45, -22, -32, -39, -35, -41, -5, 4, -26, -25, 4, 0, 12, 90, 75, -2, -8, 9, 4, 14, -35, 16, 25, 18, -14, 28, -3, 4, -5, -22, -48, -10, -38, -39, -4, -5, -33, -14, -27, -34, 4, 73, 85, 20, 9, 13, 22, 13, -24, 17, 14, 32, 26, -10, 16, -5, -17, -46, 0, 0, -34, -21, 8, 7, 10, 3, -14, -50, -38, 53, -11, -27, 17, 12, 47, 42, -8, 13, 36, 84, 29, 20, -7, 4, 6, -22, 0, 0, -45, -50, 13, 13, -2, 7, -2, 2, -44, 39, -13, -20, 0, 40, -2, 29, 8, 20, 41, 43, 23, 10, -5, -27, -6, -29, -45, -71, -82, -62, -28, 5, 33, -16, -2, -27, 3, 50, 0, 42, 24, -1, 24, 12, 1, 9, 19, 9, 12, -7, -31, -63, -19, -60, -71, -47, -72, -89, -36, -8, -20, -2, -5, -4, -9, 51, 34, 38, -19, 18, 42, 44, 1, 0, 28, 26, -17, -37, -39, -63, -54, -70, -8, -40, -82, -62, -12, 20, 6, 37, 55, 4, 25, 39, 32, 49, -5, 26, 57, 42, 9, 4, -16, -32, -9, -58, -69, -65, -30, 7, 41, -7, -61, -58, -29, 36, 25, 67, 88, 45, 2, 7, -11, 15, -16, -1, 61, 71, 11, -33, -21, -4, -42, -51, -26, -39, -26, 22, 73, 20, -11, -51, -8, 50, 71, 69, 48, -18, -24, 3, -27, 0, -3, 30, 82, 73, 40, -23, -45, -32, -30, -51, -25, -9, -16, 29, 52, 44, -12, 38, 70, 88, 67, 29, 11, -84, -59, -4, -6, -19, 8, 6, 43, 92, 47, -93, -94, -76, -42, -7, -27, 1, -33, 7, 49, 59, 42, 60, 57, 60, -4, -35, -133, -133, -136, -29, -52, -27, -12, 15, 31, 40, -61, -93, -91, -93, -3, -2, -27, -10, -53, 15, 41, 47, 22, 30, -18, -64, -105, -178, -181, -199, -111, -39, -26, -28, 19, 28, 19, -20, -143, -168, -85, -38, -37, 10, -5, 30, 25, 7, 28, 2, -50, -65, -125, -196, -222, -207, -169, -129, -68, 9, 28, -23, -7, -27, -12, -39, -149, -148, -91, -67, -50, 28, 56, 53, 49, 26, 28, -58, -103, -194, -180, -159, -151, -107, -97, -44, 23, 31, 14, -50, 14, -9, 10, -46, -135, -173, -91, -58, -30, 33, 56, 33, 28, 19, -25, -16, -28, -116, -40, -68, -97, -39, -20, -19, 89, 70, -18, 33, -48, -13, -47, -18, -91, -153, -122, -74, 1, 21, -4, -9, -16, 11, -23, 29, 21, -2, -6, -19, -38, 13, 27, 1, 104, 47, -21, 55, -17, -16, -58, -28, -117, -152, -91, -18, -15, -14, 26, 7, 6, 15, 0, 54, 35, 57, 12, -10, -6, 28, 60, 34, 31, 66, 12, 45, -6, -32, -5, -45, -123, -173, -112, -60, -42, -12, -33, -7, 36, 30, 24, 57, 37, 37, 21, 35, 28, 52, 30, 39, 55, 30, 24, 6, -6, 2, 23, -55, -115, -147, -80, -109, -66, -45, 14, -15, 25, 47, 33, 86, 93, 58, 91, 70, 63, 40, 28, 49, 1, 30, 38, 10, 15, 4, -38, -6, -29, -103, -93, -87, -49, -46, -31, -7, 33, 44, 71, 104, 87, 85, 98, 79, 73, 38, 29, -3, -57, -2, 39, -5, 18, 1, -15, 7, 8, -4, -91, -84, -95, -63, -16, 4, 42, 28, 24, -5, 14, 34, 24, 21, 12, -42, -23, -15, -13, -5, -14, 13, 16, 16, -19, -18, 13, -9, -17, -61, -63, -40, -45, -21, 29, 39, 16, -35, -32, -15, -23, -37, -43, -40, -21, -14, 12, -2, 17, -1, 7, 3, 17, 1, 7, 13, -20, -16, -13, -19, -20, 12, 3, 6, 23, 0, 10, -13, -9, -5, 20, 18, 15, 12, 18, -15, 19, 6, -16, -752, 19, -4, -12, -5, -15, 3, 18, 9, 3, 18, 28, -15, 0, 3, -23, -39, -22, -26, -17, 6, 23, -22, -5, 0, 1, 8, -5, -6, 7, -14, 13, 11, 3, -43, -37, 12, 24, 14, 8, -31, -94, -91, -110, -120, -126, -122, -77, -45, -44, -36, -19, 22, -13, -19, -9, -19, -18, -16, 15, 11, -5, -12, -32, -29, 11, -21, -74, -105, -145, -78, -78, -71, -165, -132, 22, 19, -28, -91, -91, -74, -13, 13, 0, -6, -1, 8, 35, 10, 23, -2, -11, -15, 13, -29, -32, -9, 12, -12, -38, -37, -76, -51, -24, -37, -10, -32, -46, -90, -31, 20, 17, 14, 10, 66, 8, 24, -8, -33, -49, -25, -9, -36, 41, 59, 26, 11, 21, -21, -32, -21, -24, -16, -13, 17, 44, -14, -44, 13, 7, -3, 2, 26, 36, 20, 31, -36, -59, -49, -46, -68, -20, -23, -12, 7, -12, -61, -84, -44, -22, -27, -6, 24, 93, -5, -5, 1, 7, 12, 12, 18, 24, 29, 25, -14, -45, -78, -85, -65, -98, -97, -54, -39, -54, -40, -63, 9, -30, -50, -17, 10, 46, -13, -21, 20, 19, 19, 29, 29, 21, 8, 10, -46, -96, -67, -90, -113, -128, -74, -109, -34, -36, 29, 40, 2, -26, 13, -25, 9, 5, -25, -83, 30, 45, -4, 49, 36, 19, 1, 2, -9, -50, -90, -56, -67, -105, -118, -123, -57, 24, 60, 19, -1, 38, -8, -22, -35, -35, -52, -69, 23, 7, 6, 46, 25, 19, -6, 18, -15, 5, -37, -26, -61, -142, -137, -86, -7, 66, 30, 16, 34, 11, 8, -22, -39, -12, 7, -24, -29, 12, -43, -40, -2, 5, -23, 39, 40, 16, -11, -31, -67, -169, -82, -15, 19, 70, 42, 27, 26, -17, -26, -15, 37, 38, 69, 41, -15, 24, 15, 0, -8, 7, 12, 14, -13, -14, -74, -99, -102, -90, -4, -23, 13, 60, 3, 36, -24, 8, -21, -33, 42, 73, 54, 13, 41, -11, -20, -8, -44, -39, -29, -57, -26, -53, -120, -153, -109, -87, 43, -9, 11, 35, 33, 24, -14, 1, 11, 24, 23, 8, 35, 25, 31, 0, -5, -11, -18, -42, -25, -30, -42, -56, -109, -107, -78, -6, 24, -16, -1, 47, 43, 14, -23, 33, 7, -7, -59, 24, 6, 15, 0, -15, -8, -43, -59, -61, -96, -109, -91, -54, -112, -92, -68, 26, 3, 9, 31, 62, 35, -36, -70, -6, -13, -40, -105, -23, 34, 29, -62, 1, 21, -35, -30, -35, -12, -40, -48, -37, -57, -54, -20, 19, 38, 29, 65, 53, 3, -106, -95, -61, -109, -84, -47, -19, 54, -1, -22, -19, -4, 3, 21, 41, 52, 28, 22, 30, 5, 17, 17, 33, 76, 95, 82, 15, -88, -156, -132, -130, -131, -127, -34, 18, 44, -15, 29, 13, 1, 27, 12, 88, 36, 38, 24, 6, 3, -11, 23, 47, 119, 88, 29, -51, -150, -186, -134, -120, -99, -67, -61, 26, 19, 5, 36, -10, -9, 2, 62, -54, -42, -20, -5, -33, -60, -11, 7, 57, 64, 64, -9, -93, -165, -220, -127, -47, -52, -30, -56, -14, 29, -2, -32, -53, -17, 7, 31, -71, -64, -41, -11, -17, -3, 24, 19, 42, 7, -3, -33, -62, -198, -201, -122, -61, -34, -31, -42, -4, 2, -13, -11, -15, -27, -9, -6, -124, -76, 0, 16, 5, 12, -6, -26, 4, -15, -26, -11, -51, -115, -159, -140, -57, -42, -19, -55, -17, 47, 9, -30, -47, 0, -12, -37, -125, -28, 19, 23, -6, 22, -27, -9, -47, -20, -63, -41, -120, -147, -138, -160, -117, -39, -13, -38, -15, 19, 14, -2, -8, -5, -13, -58, -104, 10, 2, 3, 0, -20, -46, -45, -37, -32, 3, -29, -99, -154, -151, -139, -137, -134, -8, -1, 25, 41, 33, 37, 10, 3, -33, -76, -74, -25, -3, -25, -36, -38, -5, -49, -48, -7, -12, -25, -80, -114, -97, -111, -108, -61, 7, 25, -3, 38, 8, 29, 12, 2, -14, -27, -45, -64, -85, -27, -56, -52, -36, -66, -82, -112, -154, -123, -132, -136, -87, -51, -35, -26, -5, 8, -21, 10, 25, 11, -20, 4, -15, -7, 15, -4, -22, -22, -14, -57, -33, -50, -84, -69, -44, -42, -56, -69, -18, -41, -47, -7, -20, -5, -2, -21, -9, 4, 19, 0, 15, -5, 11, 3, 16, 21, 12, -9, -3, -2, -83, -38, 2, 22, -5, -24, -17, -31, -18, -26, 1, -14, 10, -2, -2, 21, -16, 15, 14, -9, -19, -17, -5, 9, 6, 7, -5, 0, -17, 16, 9, -18, -14, 12, -4, 16, 9, 10, 4, 8, 15, 2, -8, -1, -7, -9, 141, 9, 4, -15, -13, 24, -11, -42, -17, -15, -16, 53, 24, -17, -17, 70, 14, 36, 17, 48, 19, -9, 4, 13, 10, 14, -12, 13, 10, 7, 10, 1, -11, -13, -52, -51, -41, 7, 3, -11, 12, -31, -51, 42, 14, 25, 38, 14, -9, -49, -88, -67, -78, 4, -17, -9, 8, 11, -6, 7, 30, -6, -54, -55, -53, 7, -5, 17, 52, 32, 15, 85, 77, 91, 89, 48, 64, 54, -6, -47, 7, -4, 12, -5, -5, 6, 28, -21, 7, -58, -75, -70, -52, -48, -17, -10, 18, 11, 43, 37, 34, 58, 41, 15, 23, 34, 15, 11, 65, 45, 27, 20, 13, 0, 29, 52, -37, -1, -38, -90, -51, -29, -1, -28, -7, -20, 0, 6, -1, 41, 29, 24, 5, 0, 14, 28, 69, 35, 80, -3, 8, -15, 23, 5, -45, -10, -28, -69, -33, -1, -25, -23, -27, -37, 2, 12, 11, -1, 4, 13, 16, -15, -47, -13, 44, -6, 3, -5, 7, -12, -7, 14, -29, 7, -27, -19, -35, 17, -22, -7, -38, -6, 39, 64, 40, 37, 13, 21, 20, 30, -21, -61, -27, 3, -20, 14, 0, 5, -21, -20, 19, 22, -4, -16, -22, -21, -6, -54, -63, -40, 18, 47, 57, 29, 37, 30, -5, 7, -10, -72, -50, 20, -9, -25, -15, -7, -30, 38, 28, 54, -20, -42, -8, -43, 0, -28, -49, -62, 47, 96, 92, 55, 34, 23, -24, -35, -5, -38, -38, -24, 13, -1, -15, -13, 26, 43, 56, 47, -30, -8, -5, 5, -21, -46, -80, -24, 42, 108, 95, 43, 17, -9, -41, -38, -20, -16, -18, 48, 32, -4, 30, -3, 3, 23, 57, 27, -41, -15, -7, -17, -55, -83, -58, 8, 77, 114, 56, 11, 11, -5, -38, -30, -28, -22, -24, 65, -14, 42, 3, -35, 31, 42, 37, 33, 2, -22, -12, -28, -39, -55, -20, 52, 112, 105, 62, 41, 25, 10, -44, -48, -40, -32, -11, 39, 1, 24, 15, -46, -11, 39, 19, 3, -21, -9, 2, -25, -48, -49, 9, 100, 128, 65, 25, 11, -24, -44, -61, -47, -26, -39, -30, 4, -5, 20, 3, 9, 17, -23, 5, 14, 6, -10, -22, -23, -44, -30, 37, 96, 73, 61, 29, -15, -21, -36, -37, -49, -40, -25, -59, 13, 59, 15, 12, -2, 104, 0, 5, -8, -40, -5, -1, -42, -7, 20, 71, 77, 105, 81, 32, 16, -40, -40, -42, -30, -11, 7, 0, 44, 50, 8, 1, 49, 84, 69, -15, -8, -38, -1, 6, -28, 22, 35, 69, 102, 110, 69, 24, 6, -15, -11, -15, -11, -29, 24, 17, 42, 58, -3, 7, 32, 79, 73, 52, 44, -15, 22, -28, -13, 22, 16, 24, 64, 94, 77, 76, 45, 1, -33, -50, -32, -32, -12, 51, 59, 99, 9, -10, 28, 62, 37, 63, 19, 13, 7, 13, -21, -8, -29, 1, 9, 46, 76, 45, 5, 9, -43, -23, -20, -45, -59, 37, 27, 30, 8, 38, 31, 81, 90, 62, 54, 68, 25, -25, -17, -23, -17, -16, -38, 13, 27, 68, 2, -30, -13, -22, -40, -20, -8, 39, 22, 12, 18, 31, 31, 27, 30, 2, 70, 58, 8, 8, 8, -27, -38, -34, -32, -13, 34, 35, 12, 3, -46, -6, -4, -24, -3, 24, 37, -27, 14, -31, 11, 45, 15, 21, 40, -15, 16, -24, -5, -12, -35, -9, -7, 8, -17, -25, -22, -23, -16, 25, 33, -27, -14, 29, 18, -12, 71, -2, 32, 69, 97, 73, 4, 6, -12, -14, -1, 39, 47, 27, 30, -13, 2, -12, -17, -13, 1, 15, 18, 22, 24, 23, 49, -19, 4, 19, 31, 52, 99, 51, 24, -24, -7, 9, 23, 17, 21, 19, 2, -32, -38, -4, -3, 3, 23, 22, 35, 2, 40, 46, 24, 42, 16, -14, 1, 51, 35, 26, -55, -65, -31, -33, -18, 42, 35, 34, -8, -28, -29, 3, 12, 38, 43, 40, 19, 20, 61, 57, 43, 12, -8, 5, 1, 12, 17, 62, 55, 44, 57, 44, 55, 26, 25, 20, 26, 9, 27, 57, 25, 54, 74, 61, 42, 63, 39, 54, 38, 4, 14, -2, -4, 18, 2, 46, 64, 48, 47, 95, 139, 130, 86, 100, 118, 66, 45, 143, 185, 145, 119, 124, 78, 43, 40, 4, 4, 5, 16, 0, 12, -5, -2, 16, 41, 46, 43, 54, 64, 78, 81, 57, 72, 0, 26, 42, 42, 54, 68, 50, 57, 57, 28, 15, 1, -7, -12, -6, 6, -7, -3, -3, 6, -21, -11, -10, -13, -18, -16, -16, 9, 14, 11, 7, -16, -3, -8, 18, -19, -4, 2, -4, -10, -5, 7, -6, 352, -11, -2, -16, -10, -33, 34, 49, 50, 69, 51, 64, 106, 108, 118, 68, 50, 56, 34, 61, 57, 17, 39, 7, 19, -2, 1, 18, -3, 8, -7, -11, 30, 8, 73, 118, 121, 135, 130, 107, 134, 134, 200, 164, 94, 97, 116, 94, 91, 116, 132, 82, 64, 9, -8, -7, -1, 17, -4, -16, 64, 78, 76, 126, 97, 96, 45, 83, 78, 52, 53, 60, 76, 21, 31, 23, 31, 42, -8, 72, 62, 22, -2, 14, 15, -18, -27, -52, 50, 88, 43, -8, -7, -30, -34, 17, -4, 7, -7, 36, 24, -16, 17, -22, -15, -9, -5, 47, 35, -55, -57, 4, -18, -3, -30, -7, 66, 76, 47, -43, -51, -84, -98, -66, -37, -22, -25, 6, -24, -25, 17, -10, 28, 8, -24, 20, 7, -30, -74, -17, -8, 7, -4, 6, 20, 67, -32, -47, -51, -98, -87, -73, -79, -50, -44, -54, -24, -41, -15, 16, 22, 9, 9, 13, -17, -41, -88, -4, 6, 14, -1, 49, 30, 15, -63, -20, -36, -63, -95, -55, -71, -59, -62, -12, -13, -26, -22, 5, -4, 3, 30, 9, 6, -77, -90, -46, 12, 29, -46, 87, 46, -18, -21, -68, -76, -67, -63, 2, -68, -48, -28, -2, -5, -39, -20, 18, 18, 0, 4, 41, -33, -128, -57, 11, 13, 0, -36, 3, 14, 12, 19, -47, -19, -48, -53, 3, -35, -17, -20, 5, -28, -41, -16, -4, 18, 44, 30, -26, 0, -135, 17, 30, 14, -28, -31, -27, -33, -28, -4, -58, -19, -26, -53, 13, -14, -21, -9, -44, -90, -32, 24, 24, 69, 40, 21, 28, -14, -85, -35, -23, 37, 25, -53, -4, 15, -15, -7, -51, -18, -64, -40, -11, -5, -37, -72, -86, -96, -30, 15, 44, 38, -11, 11, 51, 8, -21, -42, -24, 8, 9, -101, -82, -11, 7, -50, -79, -25, -46, -34, -8, -17, -75, -109, -82, -76, 3, 24, -3, 20, -16, 3, 44, -3, -27, -77, -8, -32, -32, -97, -49, 24, -6, -47, -31, 8, -15, 2, -30, -51, -57, -50, -79, -28, -18, -8, -15, -14, 34, 1, 27, -2, -30, -52, 3, 17, -38, -38, -20, 32, 12, 22, 6, 1, -11, -15, -69, -53, -34, -12, -13, -49, -49, 13, 17, 0, 12, -8, 13, 27, 25, 36, 23, 26, -57, -20, -2, -25, 26, 28, -1, -5, -22, -79, -64, -86, -64, 12, -15, -10, -3, -4, -11, -1, 3, 28, 22, 108, 46, 35, 18, 17, 24, 61, 38, 12, 74, 40, 21, 3, -2, -9, -34, -88, -4, 8, -29, -8, 25, -1, 4, -4, 24, 31, 14, 73, 39, 31, 3, 3, 56, 97, 81, 117, 111, 84, 69, 78, 22, 16, -29, -13, 37, 64, 72, 20, 42, -1, -43, 14, 25, 41, -14, 18, 5, 46, 44, 7, 52, 69, 92, 132, 81, 44, 36, 40, 41, 39, 23, 73, 99, 106, 104, 52, 34, 10, 1, -8, 2, 11, -1, -9, -47, 40, 24, 4, 15, 36, 90, 100, 72, 56, 17, 37, 46, 99, 103, 112, 90, 98, 87, 34, -21, -24, -31, -21, 28, 14, -23, -90, -16, -32, 37, 31, 37, -5, 27, 43, 23, 33, 43, 45, 76, 121, 134, 123, 70, 77, 47, 45, -13, -52, -28, -17, -9, -44, -69, -71, -39, -13, 30, 23, -2, -34, 26, -24, -18, 22, 62, 76, 45, 74, 95, 77, 73, 38, 13, -25, -68, -78, -76, -75, -63, -73, -54, -70, 6, 16, -19, 18, -1, -5, -11, -90, -81, -22, 44, 37, 31, 9, 6, -45, -46, -31, -67, -89, -66, -94, -115, -158, -106, -31, -11, -7, 38, 13, -25, 13, -38, -10, -34, -75, -96, -60, -61, -59, -89, -105, -126, -131, -116, -66, -53, -69, -83, -116, -140, -158, -152, -93, -21, -25, 0, -23, -12, -10, -8, 6, -21, -29, -36, -65, -69, -82, -53, -20, -53, -67, -22, -54, -61, -98, -98, -178, -165, -141, -123, -93, -38, -26, 47, 8, -13, 0, 2, -11, -10, -36, -62, -43, -67, -79, -98, -70, -80, -97, -54, -54, -65, -56, -78, -112, -61, -80, -50, -64, -54, 2, 8, 16, 12, -15, -8, 6, -5, -42, -23, -71, -86, -51, -53, -30, -81, -52, -142, -106, -36, -18, -35, -51, -48, -33, 0, -19, -14, 28, 1, 7, -16, -3, 13, 18, -10, -7, 23, 41, 26, 32, 25, -1, 29, 2, 22, -27, 0, 8, -4, -21, 0, 8, -11, -8, -10, 12, 17, 17, -18, 19, 6, -15, 8, 20, -17, 0, -18, 15, 16, 14, -10, 1, 5, 21, -13, -5, 2, 0, -9, -15, 10, -9, 4, 0, -16, 3, 8, 19, -1108, 11, -7, -19, 2, -14, -4, -8, -23, 18, 16, -9, -4, 49, 61, 28, 39, 34, 3, -18, -5, 12, 20, -44, 0, 4, 13, -11, -14, -20, -16, -11, -11, 5, -36, 1, 3, 12, 12, 44, 12, 18, 77, -9, 34, 20, 39, 47, 34, 82, 89, 111, 78, 22, -15, -17, -2, -13, -16, -11, 39, 56, 10, -17, -9, -18, -11, -14, -15, -53, -8, -10, -4, -21, -13, 16, -1, -4, -28, 36, 11, 37, -17, -1, 12, 21, -3, 0, 32, 35, 21, 20, -22, -41, -10, -21, -63, -78, -83, -83, -52, -44, -13, -32, 21, 17, -17, 8, -18, -65, -36, -12, -8, -20, 32, 7, 37, 5, -7, 7, 0, -18, -31, -20, -57, -97, -65, -49, -47, -31, 6, 20, 6, -11, -6, -1, -70, -70, -41, 11, -14, -18, 14, -25, 46, -1, -25, -3, -14, -45, -35, -76, -94, -65, -46, -84, -58, -31, 0, 28, 20, -26, -43, -55, -44, -58, -15, -7, 9, 3, -19, 35, 47, 22, -15, -2, -17, -80, -45, -118, -87, -82, -38, -51, -40, -21, -9, -16, -15, -56, -145, -78, -82, -50, -13, -24, 6, 29, 8, 19, 41, 11, 46, -34, -62, -71, -97, -101, -80, -60, -25, 1, 7, -34, -46, -83, -90, -123, -115, -68, -60, -46, -1, 5, -4, 16, 13, 13, -12, -47, -17, -4, -68, -88, -126, -140, -121, -69, 13, 39, 6, -40, -75, -110, -144, -170, -136, -89, -50, -19, -30, -48, 18, 16, 54, 11, -42, -12, 10, 12, -84, -118, -153, -138, -100, -2, 56, 51, 2, -21, -64, -118, -157, -177, -163, -71, -38, -28, -42, 20, 13, -71, 21, -18, -38, -4, -2, 27, -59, -122, -144, -102, 0, 13, 35, 24, 8, -4, -8, -58, -106, -172, -154, -104, -46, -29, -19, -1, -8, -60, -47, -95, -113, -85, -57, -29, -104, -161, -117, 18, 47, 10, 34, 38, 61, 48, 55, -22, -29, -100, -137, -63, -16, -56, -45, -14, 15, -31, -58, -58, -114, -87, -93, -87, -160, -127, 7, 26, 64, 41, 36, 57, 50, 57, 39, 27, -21, -86, -123, -90, -11, -35, -45, 1, -14, -10, -52, -60, -117, -137, -115, -113, -96, -67, 12, 12, 50, 51, 71, 57, 38, 4, 26, 27, 12, -20, -52, -80, -1, -29, -47, -19, -26, -30, -85, -52, -84, -123, -104, -63, -73, -34, 1, 5, 61, 67, 83, 68, -15, -37, 12, 28, 42, 42, -21, -95, -37, -37, -44, -2, -8, 12, -70, -75, -58, -55, -107, -42, -36, -26, 7, 2, 29, 55, 69, 35, -46, -42, -21, 4, 8, -29, -62, -111, -50, -54, -35, -17, -20, -8, -72, -53, -19, -22, -37, 1, 1, -23, 0, -8, 12, 52, 40, 9, -38, 2, 19, -9, 15, -64, -105, -72, -49, -60, -26, -45, -19, 6, -44, 15, 4, -2, -59, -32, -55, -24, -44, -52, -15, 43, 21, -7, -32, 10, -5, -5, -20, -104, -164, -72, -59, -39, -8, 12, -36, 12, 6, -35, 3, -39, -22, -32, -72, -59, -74, -44, -2, 26, 13, 14, -24, -15, 10, -28, -36, -108, -141, -74, -57, -48, -50, -35, -23, -42, 2, 48, 0, 3, 7, -13, -67, -30, -38, -5, 8, 32, 2, 16, 7, 5, -30, -71, -50, -101, -86, -71, -38, -37, -60, -52, -38, 10, 19, -6, -19, 6, -15, 11, 11, 38, -6, 51, 54, 36, 58, 66, 17, -23, -64, -70, -94, -131, -133, -54, -52, -43, -60, -63, -19, -13, 31, -40, -29, -57, -42, 2, -13, -18, 35, 36, 32, 19, 35, 2, -10, -46, -85, -74, -70, -113, -128, -72, -5, -18, -28, -31, -10, -26, -63, -69, -81, -59, -74, -45, -40, -13, -47, -57, -75, -71, -47, -59, -46, -49, -89, -82, -47, -33, -59, -19, 28, 22, 20, 9, 6, -47, -37, -108, -67, -41, -57, -37, -56, -8, -39, -40, -60, -71, -52, -35, -88, -79, -85, -88, -54, -23, -2, -20, 36, 32, 18, -17, 0, -4, -44, -67, -40, -89, -80, -65, -45, -56, -71, -69, -147, -145, -136, -135, -119, -127, -92, -77, -33, -15, -11, -22, -19, 17, 27, 15, 1, -20, -3, -16, -42, -16, -41, -53, -27, -21, -94, -59, -88, -85, -90, -83, -78, -71, -102, -52, -40, 9, 9, -9, -17, -21, -19, -16, -1, -3, 18, 14, -20, -27, -3, -4, -21, -44, -15, -42, -45, -46, -21, -16, -8, -32, -20, -24, 3, -28, -7, 0, 0, -7, -2, 11, 14, -17, 0, 18, -4, -1, -13, -5, -3, 0, 7, 9, -15, 13, 2, -1, -1, 19, 20, -6, -7, -7, 9, 18, 0, -6, 2, 5, 0, -999, 0, 10, 0, 13, 1, -10, -7, 1, 19, 36, 1, -6, -21, -53, -19, -5, -8, -23, -18, -5, -24, -4, 13, -15, 6, 5, -7, -8, -8, 13, 9, -3, 15, -4, -37, 5, 13, -4, -3, -41, -86, -103, -100, -99, -90, -82, -42, -39, -52, -22, -17, -13, -15, -7, -14, -9, 9, 13, 10, 10, 27, 6, -16, -20, -15, 7, -28, -60, -115, -87, -27, -70, -110, -78, 18, -8, -55, -88, -96, -62, -20, 19, 4, -9, 15, 22, 28, 9, 28, 21, -3, 5, 15, 29, 38, 2, -21, -39, -30, -8, -34, -64, 13, -46, -21, -19, -22, -77, -32, 7, 15, 18, -18, 66, 48, 39, -2, -24, -39, -4, -27, 5, 58, 25, -9, -16, -6, 12, -32, 9, 0, 17, 5, 66, 73, -16, -4, -9, -5, 3, -15, 20, 23, 19, 7, -47, -42, -47, -27, -51, -27, -2, -36, 0, -9, -51, -89, -48, 15, -13, 20, 44, 87, 30, -1, -4, 5, 23, 17, 33, 24, 24, 24, -29, -72, -50, -55, -83, -70, -58, -57, -35, -63, -59, -45, -4, 1, -13, 2, 31, 81, 20, 3, -15, 23, 6, 12, 6, 10, 14, 14, -49, -60, -83, -51, -69, -109, -70, -93, -66, -51, -13, 14, -27, -32, 14, 5, 4, -1, -3, -32, -6, 5, 0, 40, -7, 9, -4, 21, -30, -46, -45, -55, -88, -70, -85, -111, -72, -22, 18, 12, -15, -15, -23, -35, -44, -68, -23, -10, 33, -6, 0, 35, 10, 24, -35, 8, 5, 26, -18, -5, -34, -110, -159, -95, -38, 15, 35, 13, -10, 8, -21, -67, -109, -110, -49, 5, 8, -8, -33, -13, -11, -10, -13, 10, 18, 6, 2, -19, -82, -166, -116, -82, 12, 21, 23, 34, 2, 5, -8, -33, -26, -41, -24, 47, 13, 14, -16, 17, -13, -11, 27, -12, 8, 10, -19, -68, -120, -133, -47, -16, 19, 55, 10, 30, 8, 32, -4, 1, -3, -3, 19, 7, 60, -8, 18, -15, -47, -49, -11, -31, -39, -32, -94, -100, -137, -97, -1, -22, 2, 25, 3, 10, -9, 40, 39, 46, -32, -30, -6, 10, 36, 7, -9, -14, -27, -6, -5, -21, -7, -17, -63, -68, -112, -42, 36, 23, 28, 33, -8, 3, -22, -14, 36, 12, -40, -28, 10, 9, 38, -15, -1, -30, -61, -73, -60, -80, -74, -16, -39, -46, -28, 0, 12, -3, 41, 37, -18, -73, -76, -21, 0, 13, -52, -54, 38, 23, -47, -5, 3, -29, -72, -62, -12, -32, -42, 25, -30, -13, -25, -4, 24, 68, 83, -2, -35, -132, -90, -71, -66, -55, -26, -15, -1, -21, -9, -16, 1, -16, -18, -24, -4, -33, -12, 11, 15, -1, 29, 14, 67, 89, 21, -18, -101, -135, -107, -87, -98, -79, -22, 17, 19, -9, 35, 12, -1, 38, -24, -13, -55, -40, -41, -15, -16, -23, -1, 26, 63, 101, -12, -92, -175, -153, -98, -54, -75, -58, -46, 12, -4, -10, -9, -1, -20, -15, -1, -111, -94, -78, -30, -22, -74, -45, -10, 43, 73, 33, -34, -101, -131, -141, -113, -53, -47, -37, -40, -31, 12, -22, -10, -15, -1, -14, -22, -129, -123, -62, -13, -33, -4, -18, 18, 59, 25, -7, -43, -114, -130, -133, -98, -65, -25, -25, -39, -16, -8, 13, -26, -17, -7, -34, -9, -137, -86, -2, 37, 8, 11, 19, 3, 11, -14, -52, -57, -92, -94, -109, -100, -68, -70, -46, -62, -20, 18, 2, -27, -23, -2, -27, -38, -92, -16, 27, 18, 11, 39, -20, -24, -38, -36, -84, -85, -98, -98, -88, -130, -108, -67, -17, -33, -8, 57, 39, 18, -18, 8, -19, -57, -113, 14, 3, 26, 17, -5, -32, -44, -36, -32, -1, -44, -105, -123, -106, -112, -113, -94, -40, -11, 13, 8, 54, 46, -10, 12, -31, -64, -99, -61, -26, -23, -14, -4, 27, -15, -50, -13, -42, -32, -60, -72, -65, -77, -85, -37, -7, 16, -9, -1, 20, 16, 16, 5, 2, -14, -41, -65, -60, -18, -61, -64, -10, -54, -90, -79, -124, -106, -82, -90, -60, -30, -34, -21, -13, -11, -24, 1, 27, 20, -9, 10, 13, 2, -13, 0, -15, 3, -7, -6, -51, -60, -59, -35, -6, -15, -29, -30, -33, -14, -15, -18, 1, 1, -22, 14, -2, 17, -13, -8, 20, -7, -6, -9, -12, 11, -5, 16, 4, -14, -41, -17, 23, 51, -27, -22, 13, 7, -17, -30, -20, 15, 14, -5, -2, 6, -3, -8, -14, -6, -4, 15, -6, -8, -5, 7, 12, 1, 0, -13, -15, -10, 0, -20, 3, 8, -1, -17, 15, -8, -10, 18, 12, 17, -11, -12, -797, -11, 7, -12, -18, -40, -49, -58, -46, -20, -53, -45, -44, -32, -43, -52, -23, -12, -40, -30, -46, -46, -48, -5, -4, -16, 15, 11, -14, -15, -18, -13, 7, -22, -59, -74, -65, -67, -88, -72, -115, -130, -108, -107, -118, -121, -123, -150, -106, -102, -106, -54, -12, 13, -1, -14, -2, -9, 22, 13, -42, -72, -68, -87, -87, -108, -94, -116, -107, -126, -94, -107, -141, -116, -117, -96, -95, -99, -95, -75, -34, -13, 21, 20, 18, 14, 11, 36, 0, -71, -12, -27, -62, -82, -10, -13, -18, 4, 12, 5, 44, 2, 10, 15, 30, 14, -26, -13, 11, 0, 7, 0, 12, -20, -12, -29, -22, -35, 0, -11, -50, -47, 7, 17, 23, -30, -2, 4, 26, 77, 84, 68, 36, 27, 17, 0, -28, 18, 49, -1, -20, 26, -11, -7, -30, -39, -13, -20, -36, 9, 8, -19, -8, -29, -31, -31, 5, -3, 35, 39, 5, 40, 36, 39, 20, 82, 48, -4, 8, -13, 24, 11, -52, -19, 3, 23, -1, -22, -48, -41, -30, -11, -37, -66, -48, -20, 21, 31, 16, 2, 19, 29, 47, 90, 67, 28, 6, -2, -18, -14, -71, -70, 10, 24, -12, -39, -41, -18, -31, -37, -69, -21, 5, -2, 23, 29, 33, 48, 27, 51, 82, 98, 35, 20, 7, 15, 21, -30, -78, -9, 35, 17, -31, -34, -48, -36, -41, -23, -44, -22, -34, -47, -14, 62, 71, 45, 10, 36, 29, 44, -21, 37, 4, 18, -5, 11, -53, 11, 21, 3, -3, -30, -31, -18, -21, -41, -28, -89, -106, -75, -4, 66, 76, 46, 20, 30, 62, 45, 17, -2, -24, 57, 32, -30, -53, 0, 27, 4, -23, -19, -2, -32, -15, -8, -30, -40, -28, -11, 9, 50, 64, 46, 36, 44, 46, 33, 39, -25, -9, 58, 98, -3, -9, -1, 9, 19, 18, -12, -15, -5, -20, -17, -37, -15, -32, -6, -9, 55, 63, 39, 40, 69, 56, 26, 31, 5, -20, 25, 78, 20, 21, 27, -6, 43, -1, 24, -29, -8, -42, -29, -15, -21, -33, -23, 9, 52, 50, 55, 29, 83, 76, 31, -6, -44, -7, 44, 74, 35, 21, 23, -2, 33, 13, 12, -32, -45, -94, -45, 0, 0, 4, 11, 32, 51, 51, 55, 53, 33, -8, -12, -38, -37, 15, 45, 50, 26, 30, 35, -5, -16, 13, 18, 15, -82, -96, -73, -26, 26, 41, 39, 28, 25, 51, 21, 27, -44, -43, -27, -43, -10, 6, 15, -44, -9, 57, 35, -4, -15, 19, -15, -37, -107, -101, -87, -35, -8, 4, -15, 14, 19, -24, -20, -31, -69, -75, -76, -58, -41, 7, -36, -65, -5, 44, 44, 41, -3, 21, -21, -56, -100, -85, -76, -31, -32, -52, -39, -59, -90, -42, -42, -41, -94, -105, -84, -65, 9, 10, -6, -38, -63, 16, 58, 74, 22, 45, -11, -22, -4, -30, -27, -53, -60, -74, -85, -83, -68, -69, -70, -75, -78, -61, -56, -22, -21, 15, -47, -109, -48, 19, 59, 49, 11, 58, 24, 5, -24, 2, -39, -39, -70, -73, -50, -55, -30, -40, -54, -36, -82, -20, 2, -4, -28, 0, -36, -119, -96, 16, 30, 32, 17, 49, 65, 22, 16, 31, 4, -38, -46, -24, -36, -21, 1, -53, -16, -5, -29, -7, 23, 2, -8, 9, 22, -138, -65, 36, 80, 78, 48, 20, 57, 70, 47, -6, -19, -42, -30, -35, 13, 24, -37, -53, -20, 0, -28, -3, 1, -17, 21, 3, -11, -110, -128, -47, 15, 95, 40, 34, 25, 44, 45, 4, -5, -39, -22, -3, -31, -37, -73, -77, -19, -10, -49, -23, 17, 17, -7, -18, -11, -46, -68, -62, -24, 53, 65, 22, 59, 74, 68, 76, 44, 6, -6, -6, -11, -51, -38, -23, -18, -16, -63, -23, -10, -4, -20, -3, 30, -58, -89, -69, -9, 9, -37, 1, -13, 23, 46, 83, 74, 33, 21, 16, -4, -25, -14, -30, -38, -45, -44, -55, -24, 20, 16, 8, 14, -17, -28, 9, -44, -53, -69, -25, -9, -9, 59, 93, 68, 98, 36, -9, 8, -19, -27, -34, -34, -24, -38, -32, 1, 3, 15, -21, -16, 4, 4, 25, -33, -29, -7, -48, -26, 4, -9, 52, 16, -15, 19, 13, -52, -43, -27, -52, -26, -10, -30, 16, 27, -20, 7, 13, 11, -20, 17, -13, -29, -60, -62, -71, -47, -52, 25, 53, 12, -11, 9, 2, -13, -6, -1, -27, -8, -23, -17, 2, 10, 18, 6, 6, 12, 4, -21, 7, 5, -12, -11, -5, 18, 3, 20, -18, -3, 8, 13, 7, 6, 12, 13, -15, -16, 10, 13, -2, 16, -7, -6, 8, -1502, 8, 12, -3, -1, 0, 6, 12, 7, -6, -6, -21, -71, -46, -89, -58, -49, 15, 8, -48, -51, -23, -45, 9, 22, -17, 5, 1, -6, 18, -16, 0, -5, -5, -31, -3, 22, -34, -44, -38, -52, 5, 19, 10, 6, 1, 2, 52, 67, 59, 80, 26, 25, 18, 14, -18, -12, 6, -3, 1, -34, 1, 31, 2, -12, -41, -29, -25, -32, -9, 1, 6, 11, 23, 4, -11, 18, -6, 4, 12, -5, 5, 15, 17, -8, 12, 5, 39, -38, 55, 32, 66, 50, -17, 5, -8, -47, -33, -37, -34, -37, -27, -4, -15, 27, 6, -4, -11, -47, -66, -28, -4, -7, 14, 17, -3, -54, -25, 16, 64, 13, -2, -9, -41, -53, -30, -32, -57, -64, -15, -12, -19, 16, -2, -34, -50, -77, -99, -67, -16, -13, 20, 54, -23, -20, -27, -11, 15, -19, -3, -31, -54, -49, -23, -68, -38, -61, -34, -18, -35, -33, -63, -93, -83, -77, -117, -80, 18, 1, -19, 31, -38, -49, -89, -65, -34, -54, -42, -62, -52, -21, -62, -43, -12, -17, -48, -82, -55, -57, -62, -98, -50, -89, -83, -85, -24, 6, 2, 7, -43, -60, -166, -122, -96, -66, -48, -31, -62, -12, -9, 15, -2, -14, -26, -94, -113, -105, -99, -57, -68, -4, -31, -14, -24, 2, 8, -38, -74, -122, -176, -154, -55, -77, -70, -28, -50, 16, 3, 31, -14, -17, -3, -82, -82, -121, -77, -55, -41, 15, 20, 2, -9, 1, 13, 33, -81, -72, -56, -87, -39, -57, -9, 20, 18, 28, 42, 50, 2, 0, 15, 17, -17, -38, -112, -91, -76, -4, -17, 49, 7, 12, -50, -24, -62, -34, -28, -68, -27, -22, -13, 52, 64, 70, 42, 36, -1, -30, 19, 42, 45, 10, -20, -85, -78, -34, -65, 29, -12, 8, -16, -41, -55, -71, -68, -65, -66, 13, 68, 68, 79, 84, 47, -2, -24, 13, 72, 44, 41, 47, 14, -81, -71, -40, -44, -12, -14, 0, -44, -22, -62, -105, -24, -26, -17, 72, 82, 85, 69, 79, 25, -30, -44, 26, 50, 66, 56, 58, 12, -56, -57, -9, 2, -8, 14, -35, -34, -102, -78, -113, -117, -56, -33, 57, 67, 61, 28, 48, 17, -36, -21, 46, 53, 92, 85, 45, -2, -78, -35, -3, 37, -12, 0, 0, -38, -78, -69, -95, -124, -84, -29, 4, 29, 30, 36, 6, 7, 4, 53, 87, 74, 80, 47, -17, -26, -62, -60, -20, 4, 1, -19, -7, -37, -80, -94, -136, -109, -100, -46, -8, 51, 39, -11, 44, 20, 44, 102, 119, 104, 55, -15, -27, -75, -72, -116, -89, -14, -16, 8, 12, -6, -120, -141, -147, -126, -82, -48, -46, 11, -9, -5, 12, 6, 26, 75, 51, 49, -31, -57, -49, -63, -87, -71, -93, -51, -27, -20, -10, -37, -59, -29, -55, -82, -92, -83, -61, -36, -61, -53, 2, 17, -9, 24, -9, -39, -57, -61, -51, -56, -44, -67, -63, -83, -37, -8, 2, 14, -50, -89, -70, -67, -62, -74, -66, -46, -37, -71, -35, 37, 35, -2, -14, -44, -44, -43, -28, -11, -48, -11, -3, -30, -39, 11, 4, -50, -30, -7, -52, -71, -24, -49, -58, -79, -35, -25, -3, 22, -1, -25, -29, -17, -11, -19, -10, -20, 9, 34, 35, -21, 42, -37, -15, 27, 52, 23, 19, 6, 13, -19, -15, -8, -5, 28, 19, 4, 8, -7, -26, -27, -35, 3, -31, -13, 17, 0, 32, -7, 33, -44, -13, 2, 2, -4, -5, -25, 9, -8, -15, -14, -1, 17, -1, 6, -6, -26, -20, -35, -35, -7, 13, -6, 28, 45, 27, -39, 0, -40, -9, 20, -26, -38, 25, 51, -36, -34, -41, -17, 19, -41, -44, -28, -31, -35, -42, -53, -22, -29, -14, -38, -41, 34, -16, -66, -27, -2, -12, -19, -49, -18, 33, 51, 53, 16, -24, -44, -49, -52, -67, -46, -59, -56, -68, -90, -114, -94, -97, -67, -9, 14, -14, -75, -10, 20, -10, -8, 18, -2, 12, 2, 47, 40, 26, -3, -30, -4, 15, 7, 9, -57, -95, -14, -40, -47, -85, -51, -20, -17, -25, -17, -33, 15, 10, -19, 4, -31, 31, 33, 54, 38, 47, 50, 6, -19, -18, 31, 45, -16, 12, 23, -4, 6, 24, -16, -30, 9, -24, -30, 10, -4, 14, -2, -14, 12, 20, -24, -25, 2, 39, 36, 37, -18, -59, -50, 16, 22, 19, -13, -9, -12, -15, -42, -30, 11, -15, 12, -11, 15, -15, -4, -7, 12, 18, 13, -6, -18, 19, -20, -1, 1, 17, -16, -12, -20, -10, -12, -12, 5, 3, 14, 21, -17, 14, -12, -14, -20, -7, -185, 15, -2, -9, 17, -21, 9, 9, 12, 57, 51, 30, 10, -29, 82, 28, 12, 30, 47, 41, 25, 24, 2, -3, -1, -8, -8, -18, -19, 9, -11, 11, 22, -27, 7, 23, 28, 25, 2, -18, -38, 32, 78, 82, 81, 35, 4, 32, 45, 39, 92, 62, 46, 15, -2, 13, 11, -15, 36, 29, -37, -65, -19, 16, 20, 20, 4, -22, -36, -5, 11, 13, 7, 38, -40, -87, -99, -75, -66, -18, -4, 38, -9, -6, 13, -20, 22, 54, 92, 30, 30, 20, -41, 16, 19, -4, -31, -17, 8, 27, 28, 11, -25, -43, -13, -39, -55, -30, -82, -80, -38, 13, 3, -5, -75, 11, 87, 26, 41, 5, -49, -27, -47, -36, -45, -54, -28, -7, 27, 39, 30, 45, 48, 17, 50, 19, -22, -83, -48, 17, -14, 3, -23, 46, 86, 28, -9, 7, -46, -57, -38, -43, -56, -32, -7, 9, 20, 25, 49, 37, 30, 42, 47, 53, 12, 9, 26, -6, -23, 15, 41, 83, 118, 62, -30, -8, -51, -42, -64, -31, -49, -41, -38, 26, 8, 33, 13, 17, 13, 2, 2, 41, 5, 6, 9, 17, -1, 13, 83, 52, 71, 42, 8, -16, -3, -40, -72, -36, -10, -29, -48, 36, 80, 78, 44, 14, 1, -4, -36, -10, -16, -66, 9, 3, -4, 18, 70, 63, 32, 42, 37, 4, -10, -49, -35, -46, -62, -83, -30, 47, 73, 57, 60, 16, 39, 27, -18, -50, -39, -67, 8, 17, -9, 12, 6, 92, 17, 32, 5, -8, -42, -45, -56, -51, -78, -57, -43, 27, 56, 41, 66, 23, 38, 18, 9, -45, -53, -93, -85, -3, 40, 69, 75, 85, -27, -59, -24, -20, -25, -63, -88, -59, -39, -16, -16, 19, 60, 52, 49, 35, 1, -1, 18, -21, -28, -59, -63, -31, 1, 69, 93, 77, -14, -25, -16, -4, -49, -70, -40, -25, -12, -40, -33, -14, 31, 41, 75, 17, 21, -12, -4, 6, -3, -63, -20, -17, -15, 45, 45, 62, 36, -30, -5, -12, 9, -37, -49, -40, -56, -31, -3, 0, 22, 32, 53, 2, -15, 15, -49, 27, 28, -36, -62, -31, -11, 41, 93, 72, 52, 22, 19, 37, 30, 0, -5, -60, -74, -40, 9, 12, 33, 39, 53, -12, -5, 0, 2, 17, 6, -40, -5, -34, -13, 40, 73, 46, 43, 25, 46, 42, 15, -28, -55, -103, -76, -69, -57, -45, 4, 0, 31, -19, -8, 6, 2, 10, 18, 7, 66, -22, 0, 45, 44, 79, 91, 69, 64, 39, -1, 0, -89, -116, -134, -83, -79, -69, -32, -34, -22, -11, -6, -2, 58, -17, -7, -25, 54, -25, -9, -4, 18, 34, 87, 92, 63, 32, 0, 1, -59, -122, -98, -68, -37, -39, -40, -9, -5, -23, 4, 10, 52, -4, -64, -16, 24, 40, 0, 21, 11, -68, 12, 39, 1, 25, 9, 39, 12, -12, -35, -9, 17, 20, 23, 33, 13, 9, -14, -32, 16, 6, -30, -12, 30, -12, 21, 24, -54, -88, 11, 48, -29, 19, 32, 80, 70, 68, 42, 54, 41, 45, 17, -13, 17, 25, -39, -56, -42, -45, -49, -7, -3, 32, 18, 14, -74, -110, 2, 29, 12, 23, 42, 55, 47, 103, 113, 38, 37, -15, 15, -17, 41, 23, -4, -58, -22, -78, -38, -25, 6, 39, 45, 20, -78, -77, -18, 29, 43, 45, 19, 27, 74, 46, 88, 27, -9, -1, 2, 3, 6, 3, -29, -60, -37, -36, -17, -58, 16, -36, 13, 7, -98, -90, -90, -42, 8, 51, 6, 27, 52, 43, 45, 50, 11, 2, -10, -10, -3, -25, -18, -23, -20, -57, -75, -61, -15, -9, -11, -35, -57, -81, -77, -86, -55, -13, -24, -13, 18, 5, 0, 3, 16, 31, 5, 17, 27, 12, -9, -19, -25, -69, -77, -55, 0, -16, 4, 14, 3, -61, -96, -43, -64, -61, -56, -77, -31, -2, -34, -25, -10, -35, -7, 29, 21, 22, -31, -47, -43, -65, -39, -16, -34, 17, 3, -17, 6, 16, -10, -3, -15, -84, -97, -80, -89, -20, -6, -43, -44, -13, 7, -9, 3, 18, -37, -27, -30, -50, -45, 23, -24, -18, -18, -3, -14, 33, 3, 20, -31, -76, -113, -108, -120, -92, -68, -53, -48, -30, 10, -22, -8, -9, -2, 30, -9, -18, -18, 2, 20, -6, 20, -13, 14, -1, 10, -10, -9, -39, -42, -61, -35, 33, 40, 42, 1, -8, 15, 32, -46, 4, -18, 16, -20, 6, -22, -20, -5, -13, 2, 7, 10, 8, -6, -8, -1, 5, -13, 10, -4, 6, -1, 22, 20, 2, 8, -16, 10, 10, -17, -15, 1, 3, -1, -15, -19, 12, -9, 1377, 2, 0, 4, 7, 0, 0, -13, 5, -28, -52, -102, -53, 4, -33, -77, -18, -5, -54, -71, -38, -44, -35, -4, -24, -19, -13, -1, 4, 12, 18, -7, 8, -4, 31, 27, -33, -27, -29, 23, 12, 26, -34, 3, 35, 18, -44, -39, -48, -63, 4, 27, 66, 26, -4, -17, -19, -4, -12, -21, 72, 75, 70, 90, 14, 18, 17, 35, 54, 28, -3, 12, 13, 56, 10, -28, -42, -40, -8, -31, -24, 11, 26, 20, 18, -17, -39, -46, 22, 58, 56, -16, -2, -11, 1, 29, -3, 20, 3, 15, 14, 9, 5, 19, 24, -5, -9, -28, -18, 14, -47, 2, -10, 5, 17, 13, 52, 39, -8, -31, 1, -31, -39, -14, 34, 8, 43, -12, 19, -1, -14, -37, 0, -24, 25, 32, 26, 5, -29, -16, -11, -6, 35, 32, 43, 33, 7, -6, -7, 4, -10, 19, 22, 23, 35, -9, 20, -7, -11, -30, -27, -23, -39, 25, 19, -43, -111, 7, 10, -1, 44, 7, 48, 10, 15, 29, 41, -10, 10, 19, 11, 36, 12, 31, 30, 29, -8, 5, -4, -25, 2, 26, 24, -74, -65, -41, 0, 11, -49, 7, 7, -9, -19, -9, -21, 22, 9, 24, 36, 7, -21, 7, 52, 46, 10, 5, -36, -51, 9, 56, -16, -55, 14, 39, 12, -25, -47, -32, 25, -3, -31, -20, -7, -18, 14, 38, -4, 3, -2, 32, 55, 100, 22, -24, 9, -10, 10, 36, 30, -16, 17, -9, 4, -21, -82, -33, 16, -16, -50, -11, -15, 20, 21, 28, 23, 9, 4, 16, 42, 42, 25, -14, 0, 11, 68, 95, 42, -57, -22, -18, -38, 6, -78, -37, -32, -8, -6, 4, 25, 48, 57, 49, -21, -14, -35, -32, -4, 6, 7, -7, -6, 35, 77, 105, 61, -6, -43, -27, 5, -56, -54, -9, 0, -25, -7, 11, 18, 39, 26, 5, -39, -47, -48, -34, -6, 43, 32, 1, 17, 12, 76, 110, 73, 2, -65, -17, -18, -25, -42, -16, 35, -23, 4, 62, 56, 56, 36, -12, -61, -95, -82, -51, 19, 19, 56, 28, 19, 79, 88, 122, 53, -32, 8, -7, 6, -54, -79, -37, 14, 4, 44, 45, 83, 36, -31, -75, -60, -67, -86, -54, 6, 44, 75, 66, 37, 76, 91, 115, 26, -27, -34, 0, 17, -30, -73, -72, -9, 50, 86, 103, 86, 22, -48, -82, -85, -82, -83, -74, 34, 37, 30, 17, 19, 36, 52, 78, 13, -36, -24, 12, 16, -55, -9, -39, 18, 115, 119, 79, 59, -14, -46, -62, -66, -64, -89, -31, 21, 61, 28, 27, 38, 58, 76, 29, -8, -38, -31, -27, -6, -52, -35, -8, 89, 101, 92, 54, -15, -33, 3, 17, 24, -54, -77, -74, 23, 8, 28, 21, 26, 27, -5, 13, -19, -60, -74, 0, -11, -57, -12, 32, 129, 82, 36, -12, -18, -44, -22, 0, -6, -20, -94, -71, 14, 7, 46, 31, 52, 27, -27, -7, 9, -94, -69, -47, 4, -48, -30, 52, 86, 90, 52, 13, -2, -43, -11, -21, -32, -41, -89, -52, -4, 24, 23, 16, 21, -6, -7, -43, -74, -59, -30, -25, -13, -9, -6, 28, 105, 120, 70, 33, -15, -42, -21, 3, -21, -7, -19, -41, -11, 37, 5, 33, 16, 4, -1, -14, -95, -37, -5, -51, 40, 9, -8, 18, 60, 123, 106, 33, -5, -11, -13, -10, 13, -14, -7, -1, -9, 46, 22, 34, 22, 32, -9, 37, -74, -66, -36, -60, -3, 4, 16, -44, 79, 121, 95, 33, 36, 34, 11, -31, -36, -41, -42, -15, 0, 29, 19, -3, -7, -11, -40, -9, -38, -113, 26, -24, 1, 33, 1, -27, 25, 79, 50, 47, -6, -9, -4, 10, -31, -40, -34, -43, -9, 14, 15, 14, -21, -42, -57, -47, -42, -46, -29, -12, 15, -4, -34, -4, 73, 110, 67, 34, 0, 5, 4, 7, -27, -35, -19, -10, -24, -15, 9, 1, -41, -35, -38, -42, -18, 18, -33, 3, -9, 1, 21, -8, 17, 28, 33, 52, 12, 29, 27, -19, -67, -54, -48, -16, -25, -2, 24, 44, 30, -5, 2, 6, 45, 23, 2, 10, -4, -12, -3, -34, -18, 53, 74, 104, 120, 88, 46, 15, -21, -19, -17, 11, 16, 16, 0, -9, 55, 86, 65, 31, 21, 14, -15, 14, 17, -18, -20, -6, -8, 42, 41, 76, 52, 58, 32, 26, -12, 14, -26, 59, 72, 35, 57, 35, 37, 57, 21, 7, -17, 17, 2, 9, -11, -11, 3, -8, 12, 17, 8, 16, -1, 6, -12, -14, 15, -14, 5, 21, -1, -10, 12, -15, 16, -5, -21, 4, -13, -1, 14, 12, 6, 522, -8, 14, 15, -18, 47, 11, -19, -22, -4, -28, 3, 11, -11, -42, 14, -27, -18, 24, 24, 18, 14, 28, 23, 6, 0, -9, -18, -19, 18, 10, 13, -27, -59, -44, -22, -57, -38, -102, -86, -23, 13, -21, -67, -115, -143, -91, -67, -51, -63, -60, -26, -39, 4, 2, -3, 11, -20, 7, 9, 9, 38, -4, -1, -10, -46, 1, 24, -9, 23, -32, -25, -62, -33, 0, -50, -72, -51, -8, -21, -5, 21, -37, -3, 15, 5, 23, 33, -30, 7, 48, 37, 7, 19, -12, 17, 4, -24, 5, -14, -6, -6, 25, -1, -14, -15, -11, 16, -21, -23, 3, -17, -7, 16, 32, -28, -30, 4, 7, 23, -6, 39, 14, -1, 0, -28, 23, -34, -23, -12, 11, 3, -16, -45, -23, 2, -15, -12, -16, 15, 9, 10, 44, -6, -3, 21, 20, 13, -15, 7, -33, -41, -28, -11, -63, -72, -50, -32, -5, -14, -48, -99, -92, -120, -79, -30, -44, 1, 11, 19, -29, -24, 0, -23, 25, -47, -53, -25, -35, -46, -47, -53, -97, -73, -65, -60, -79, -84, -100, -133, -176, -131, -63, -83, -64, 11, -10, 18, -16, -76, -60, -62, -73, -29, -77, -41, -52, -37, -35, -34, -60, -58, -94, -93, -108, -78, -99, -80, -53, -109, -90, -54, -2, -25, -18, 19, -34, -107, -71, -86, -107, -43, -46, -39, -38, -20, -28, -7, -3, -54, -63, -37, -62, -54, -49, -42, -23, -53, -30, 13, 4, -9, 0, -2, -47, -81, -47, -44, -64, -20, 20, -35, -34, -22, -15, 14, 55, 4, 36, -22, -26, -5, 8, 34, -10, -22, -39, -17, 46, -5, -44, -33, -52, -52, -59, 18, -21, 42, 14, 32, 57, 9, 25, 65, 54, 26, 14, 17, 6, 34, 53, 31, 25, 9, -20, -29, 0, -1, -19, -55, -51, -53, -40, -20, 12, 47, 27, 25, 19, 45, 21, 55, -18, 0, 15, 33, 12, 21, 64, 58, 24, 23, -13, 9, -14, 2, -3, -25, -11, -12, -39, -16, 29, 4, -34, -6, 0, 40, 42, 14, -31, -61, 5, 24, 25, 52, 32, 26, 37, 37, 21, 38, 38, 35, 30, -10, -54, 6, -3, -21, -7, 11, -11, 2, 18, 39, 36, 5, -34, -60, 52, 70, 25, 30, 39, 31, 47, 70, 48, -33, 45, 46, 20, -56, -26, 25, -50, -100, -24, -8, -6, -14, 3, 32, 28, -28, -61, -38, 69, 94, 46, 50, 61, 44, 24, 29, 4, -56, 24, 22, 1, -54, 33, 32, -39, -91, -13, -9, -4, -1, -7, -9, 14, 25, -33, 38, 106, 93, 73, 72, 56, 41, -6, -20, -28, -64, 18, 42, 28, -49, 8, 47, -22, -2, 2, 5, -12, -25, -22, -10, 62, 76, 19, 42, 132, 79, 89, 77, 59, -5, -44, -32, -26, -45, 70, 6, 16, -3, 5, 87, 58, 63, 80, 58, -5, 16, 18, 47, 95, 118, 81, 73, 82, 40, 52, 33, 12, 4, -17, 28, 30, -29, 57, 58, 29, 35, -12, 26, 64, 45, 58, 52, 48, 40, 41, 41, 66, 78, 17, 35, 41, 46, -5, -19, -33, 8, 11, 38, 31, -21, 55, 67, 15, -30, -64, 65, 88, 70, 63, 32, 24, -5, 17, -12, -38, -29, -72, -52, -61, -35, -11, 3, -12, 4, 29, 13, 33, 14, 87, -11, -32, -42, 27, 59, 101, 59, 26, -9, -16, -40, -75, -82, -117, -111, -110, -74, -91, -38, -52, -36, -21, -22, -6, 39, 23, 7, 15, 26, 15, -15, -15, 15, 42, 38, -8, -78, -101, -95, -112, -118, -116, -126, -87, -98, -78, -91, -119, -58, -65, -52, -43, 43, 19, -19, -20, -1, 7, -37, -90, -38, -5, -6, -31, -112, -108, -103, -77, -31, -20, -2, -13, -93, -59, -65, -74, -51, -62, -81, -78, 15, 2, 10, -53, 10, 6, -42, -52, -23, 41, -26, 1, 19, -19, -39, -64, -54, -69, -72, -70, -19, -38, -91, -122, -111, -97, -100, -99, -52, -15, -55, 0, -17, 19, 4, -24, -82, -79, -84, 16, -8, -42, -74, -71, -97, -105, -114, -95, -167, -156, -92, -131, -158, -130, -84, -76, -35, -28, -47, 3, 12, 9, -20, 20, -60, -78, -76, -41, -98, -106, -138, -93, -56, -76, -101, -68, -50, -91, -163, -74, -99, -120, -59, -54, -28, -33, 0, -15, 10, 0, 16, -18, -2, -15, -39, -38, -51, -95, -46, -92, -126, -95, -104, -32, -79, -95, -76, -70, -74, -32, -41, -68, -23, -13, -7, -15, 4, -2, -1, 0, 16, 10, 3, 9, 12, 16, 16, -3, 10, 6, 1, -14, -23, -31, -1, 14, 9, 18, -6, -6, 0, -4, 0, 7, 11, -8, -1738, -6, 14, -12, 0, 30, 12, 31, 18, 27, 40, 70, 12, 21, 46, 40, 8, 34, 44, 21, 21, 28, 13, -7, -7, -16, -9, 15, -10, -9, -6, -6, -9, 21, -15, 10, 8, 37, 64, 57, 30, -8, 44, 20, 15, 31, 61, 20, 27, 3, -11, -2, -4, 0, -20, -4, -6, -18, 23, 32, -77, -87, -75, -65, -26, -21, -11, 7, -7, -52, -8, -5, -23, -57, -18, -8, 37, 44, 94, 50, 53, -30, 13, 12, 13, -5, 12, 69, -19, -58, -45, -4, -40, 2, 1, 39, -5, -8, -4, -12, -23, -14, -35, -33, -19, 2, 18, 54, 103, 13, 24, -20, -3, -17, -12, -42, -38, -57, -25, 19, -19, 20, 17, -4, -7, -10, -28, -4, -23, -1, -19, -15, -23, -5, -52, -7, 16, 61, 47, 7, 9, -10, -13, -8, -31, -68, -11, 27, -11, 7, -32, -47, -31, -30, -12, -26, -18, -23, -33, -34, -34, -36, -30, -12, 15, 85, 53, -9, 9, 0, -32, 18, -31, -2, -11, -16, 6, 6, -7, -45, -3, -12, -38, -15, -23, -35, 14, -7, -13, -40, -56, -48, -42, 42, 24, 27, -9, 4, 27, 26, -4, -2, 7, 26, 32, 19, 11, -25, -16, -38, -13, -6, -35, -43, -1, -13, -30, 15, -54, -62, -39, 13, -13, -38, -16, 18, 60, 23, -18, -7, 41, 25, 47, 47, -2, 15, 7, -33, -10, 7, -48, -64, -7, -17, -23, -20, -59, -47, -38, -11, -9, -4, 7, 19, 69, 36, -3, 27, 33, 39, 45, 30, 19, 16, 2, -28, -13, -7, -43, -37, -16, -7, -17, -26, -30, -30, -17, 37, 67, -4, 51, 10, 96, 68, 34, 20, 20, 58, 24, 40, 1, -8, -17, -2, -5, 10, 1, -45, -32, -23, -20, -16, -24, -97, -18, 29, 39, 31, 0, 10, 86, 14, 64, 49, 39, 42, 37, 1, -18, -22, 11, -3, 6, 17, -35, -22, -16, 5, 3, -16, -47, -102, -46, 43, 29, 51, 21, 32, 77, 40, 53, 51, 35, 5, -11, -5, -41, -3, 33, 30, 1, 7, -38, -32, -41, -18, -33, -62, -24, -87, -66, 20, -7, 13, -24, 48, 96, 99, 49, 53, -26, -27, -64, -33, -18, 5, 27, -1, 12, -5, -31, -29, -40, 2, -26, -56, -108, -97, -52, -13, 21, 27, -28, 31, 95, 134, 91, -6, -57, -69, -109, -68, 1, 14, 20, 16, 57, 18, -8, -28, -4, -8, 13, -53, -53, -65, -36, -41, 63, -11, -15, 24, 43, 118, 22, -74, -103, -115, -92, -103, -22, 14, 39, 35, 71, 13, -4, -11, 0, 4, -1, -52, -95, -41, -42, 28, 36, 35, -19, 6, 29, 22, -53, -90, -132, -172, -108, -116, -29, -1, 25, 60, 68, 36, 14, 27, 9, 10, -34, -36, -4, 1, -19, 79, 43, 0, 10, 75, 5, -2, -114, -139, -154, -132, -167, -126, -37, 35, 77, 95, 104, 71, 23, 30, 17, -4, -37, -12, 19, 26, 26, 100, 41, 7, 20, 11, 23, -53, -118, -163, -158, -169, -179, -88, -25, 55, 87, 135, 108, 87, 20, -2, 19, -3, -17, -23, -11, 64, 54, 64, 62, 30, 19, 10, -11, -66, -169, -183, -191, -210, -149, -72, -34, 54, 69, 86, 63, 63, 8, -32, 4, -24, -30, -10, -5, -7, 82, 55, 25, 44, -31, -22, -38, -34, -122, -167, -209, -165, -157, -91, -36, -6, 5, 9, 10, 24, 22, -7, 12, -3, -7, -31, -9, -14, 65, 71, 26, 67, 10, 7, -50, -41, -99, -114, -178, -143, -159, -128, -38, -14, -1, 20, 27, 19, 14, 9, 34, 24, -18, -7, 34, -11, 58, 73, 6, 7, 15, -13, -31, -23, -68, -138, -161, -121, -140, -103, -60, -73, -10, 1, -6, 12, 18, 34, -9, 12, 37, 33, 36, 54, 65, 42, 10, 5, 5, -15, -6, 7, -31, -83, -116, -93, -132, -101, -103, -100, -15, -21, -18, 30, 40, -7, 25, 24, 42, 12, 44, 50, 42, 22, 49, 21, -18, -9, -33, 9, 22, -39, -89, -80, -100, -96, -113, -31, 14, 33, 35, 38, 61, 16, 19, 30, 15, 27, 17, -3, -12, 14, 9, -7, -9, -1, -15, 19, 35, 16, -45, -39, -96, -112, -102, -84, -57, -46, -11, -11, 8, -8, 4, 7, -4, -60, -46, -53, -16, -14, -17, 9, -4, -15, -12, -1, 20, -22, -19, -53, -53, -51, -41, -29, -33, -28, -5, -67, -52, -45, -54, -30, -36, -54, -57, 7, 8, 20, 10, 12, -8, -16, -13, -11, 15, -12, -14, 11, 18, -13, 10, -16, -11, 8, -10, 2, -24, -12, -21, -7, -17, 9, 17, -16, -16, -19, -20, -16, -15, 149, -11, -13, 8, -17, -7, -19, -15, -29, -12, -14, -47, -4, 5, -15, -84, -50, -41, -46, -53, -63, -19, -12, -16, -16, 10, 0, -19, 3, -19, 0, -3, 13, 33, 20, 26, -21, -18, 34, 31, -22, -12, -40, -48, -16, 13, 21, 6, -32, -17, 37, 35, 49, 8, 2, 9, -1, -4, -23, -13, -26, 20, 43, 15, 15, -10, 11, 11, -10, -36, -60, -32, -11, -17, 33, 24, -4, -10, 10, -29, -60, -30, 19, 12, -16, 12, -45, -41, -42, -14, -24, -82, -61, -69, -73, -58, 25, 8, -11, 30, 38, -8, 15, 37, 25, 16, 8, 11, 2, 68, 1, 7, -8, 4, -38, -45, -33, -51, -85, -109, -106, -155, -132, -62, -21, -6, -26, -15, -13, 11, -5, -13, -1, -7, -9, 35, 38, 69, 21, -15, 11, -14, -19, -18, -50, -44, -74, -100, -166, -206, -127, -50, -19, -36, -11, 9, -5, 43, -7, 15, -27, -4, 1, -10, 16, 2, -33, 15, 22, 16, -18, -29, -72, -90, -103, -125, -134, -151, -71, 35, -15, 10, -27, -11, -8, 15, 33, 5, 18, 26, 57, 26, 19, -2, -54, -24, 3, 31, -25, -36, -80, -79, -97, -153, -149, -97, 8, 81, 22, -25, -7, -31, -40, -29, 15, -3, 41, 31, 67, 50, 33, 21, -25, 36, 11, -1, -14, -5, -42, -88, -149, -151, -109, -56, 53, 77, 39, 14, 6, -34, -67, -72, -11, 4, 59, 27, 53, 61, 7, 27, -13, -19, 16, -30, -15, -38, -80, -130, -136, -125, -91, -16, 61, 89, 59, 16, -10, -51, -100, -59, -55, -46, 31, 57, 85, 78, 54, 49, -6, 31, -44, 11, -53, -61, -90, -81, -106, -53, -24, 12, 62, 49, 16, -9, -69, -97, -107, -128, -146, -101, -52, 18, 32, 53, 93, 65, -6, 39, -2, -6, -69, -52, -72, -76, -84, -56, -12, -8, 33, 11, -38, -41, -22, -41, -59, -98, -140, -149, -128, -70, -28, 11, 40, 6, 38, 45, -7, -36, -89, -83, -65, -66, -26, -53, -6, -24, -2, -35, -21, -33, 15, 38, 19, -43, -87, -126, -133, -111, -76, -83, 11, -21, 40, 21, -14, -14, -75, -98, -99, -122, -53, -45, -10, -46, -41, -23, -6, -13, 20, 72, 14, -27, -71, -98, -72, -83, -107, -93, -54, -34, -55, 15, 5, -37, -60, -90, -128, -144, -120, -73, -13, -26, 5, 6, 2, 46, 65, 61, 44, -22, -22, -64, -34, -51, -54, -126, -53, -26, -65, -24, 23, -40, 20, -11, -94, -66, -118, -73, 11, 4, 41, 44, 24, 49, 82, 75, -6, -15, -11, -41, -13, -51, -43, -111, -77, -97, -66, -24, 2, -28, 48, 92, 68, 2, -23, -41, -9, 10, 67, 52, 43, 77, 70, 32, 2, -40, -38, 2, 4, -13, -58, -127, -80, -85, -97, -7, -28, -21, 43, 51, 98, 61, 6, -10, 1, -14, 32, 11, 27, 9, 38, -34, -21, -8, -19, 35, 22, -30, -99, -113, -47, -49, -55, -12, -13, 2, 57, 79, 69, 14, 8, 10, 3, -6, -16, -4, 4, -30, -44, -39, -40, -13, 33, 17, 11, -58, -51, -86, -35, -28, -2, -53, -20, 32, 67, 90, 51, 19, -6, -6, 2, -34, 10, -7, 6, 13, -4, -12, -19, 7, 2, -13, -66, -54, -35, -23, -32, -22, -59, -54, -14, -7, -1, 18, 26, 25, -18, -19, 8, 1, 8, 16, 30, 27, 2, -11, -6, -2, -48, -70, -74, -104, -115, -34, -36, -40, -24, -43, -18, 13, 28, 42, 55, 25, 2, -34, 18, 1, -19, 2, -10, 1, -2, 25, -22, -27, -81, -90, -94, -113, -126, -67, -62, -49, 4, 13, -9, -7, 59, 22, 3, -2, 39, 32, 33, 4, 12, 39, -19, 5, 9, 1, -42, -38, -71, -116, -138, -74, -54, -42, -29, 53, 0, -1, -11, 21, 56, 5, 36, 11, 18, 32, -1, -19, -7, 4, -16, 32, 21, 12, -22, -31, -96, -99, -85, -44, -31, 14, 2, 8, -14, -8, 19, 19, -15, -12, -6, -14, 8, 29, 44, 8, 16, -15, -37, 14, 19, -8, -29, -49, -62, -40, -34, -10, -14, 19, 44, 7, -33, 3, -9, 18, -19, -22, -41, -52, -19, -25, 0, 13, -15, -19, -31, -49, -74, -42, -32, -63, -66, -62, -27, -25, -10, 10, 19, 5, -7, 3, 0, -2, -6, -5, 12, -8, 0, 32, 19, 18, 11, -58, -50, 32, -9, -21, 9, -16, -18, 3, -17, 0, 18, 4, -3, 13, -8, 13, -16, 8, 16, 4, 6, -15, 14, -8, -17, 7, -7, -5, -16, 3, -16, 3, 4, 11, -2, -14, -18, 12, -3, 11, -18, -12, -16, 10, -20, 661, -5, 15, -16, 1, 26, 20, 39, 29, 65, 36, 85, 63, 71, 44, 92, 21, 43, 38, 32, 23, 10, 18, -4, 9, 6, 5, -3, 13, -2, -19, -6, -18, -36, 3, 13, 38, 55, 46, 92, 79, 93, 99, 36, -12, -4, 6, 38, 33, -1, 5, -3, -33, -5, -11, -5, 4, 12, -8, 29, 5, 55, 45, 30, 21, -19, -3, -11, -33, -22, -30, -57, -36, 1, -25, -26, -27, -70, -38, 22, 44, 26, -10, -1, 3, -7, -7, -8, 10, 61, 44, 98, 14, 8, -17, -39, -65, -70, -52, -59, -77, -37, -33, -36, -29, -56, -8, 38, -26, -58, -41, 1, -14, 0, 19, -4, 25, 37, 5, 25, 23, 9, -1, -15, -39, -37, -6, -40, -10, -42, -36, -47, -81, -18, 14, -6, -39, -88, -51, -9, -8, -2, 6, 17, 76, 14, -3, 17, -19, 9, -44, -37, -49, -55, -69, -44, -55, -66, -54, -89, -74, -77, -32, -13, -40, -73, -47, -20, 15, 8, -43, 14, 115, -4, -54, -29, -57, -37, -75, -71, -55, -85, -90, -126, -106, -136, -103, -124, -147, -129, -83, -37, -32, -65, -17, -29, 18, -21, 16, 40, 36, -47, -72, -65, -57, -66, -49, -59, -29, -67, -81, -74, -73, -78, -63, -90, -86, -88, -98, -71, -23, -51, -32, -53, -8, 14, 35, 7, -19, -69, -79, -28, -12, -7, -55, -70, -70, 16, 18, 9, 11, 35, -17, -9, 20, 14, -58, -1, -1, 20, -22, 5, 4, 43, 76, 36, -40, -20, -22, -19, 1, -6, -41, -34, -11, 73, 95, 80, 82, 86, 79, 78, 49, 23, -11, 35, 17, -52, 23, -1, 5, -33, 77, 45, 30, 30, 13, 18, 12, 5, 21, 17, 37, 68, 62, 36, 88, 39, 54, 65, 79, 70, 41, 26, 21, -48, 23, -14, -7, 3, -9, -38, -38, -17, -29, 20, 8, -27, 24, 45, 51, 29, 3, -18, 13, -25, -12, 13, 80, 98, 62, 36, 21, -18, -13, -36, -2, 51, 84, -9, -19, -16, 6, -17, -33, -25, 22, 86, 50, 18, -18, -12, -41, -36, -4, 8, 59, 76, 77, 32, 53, 79, 27, 3, 3, -7, 28, 9, -33, -12, 2, 2, -14, 36, 77, 70, 30, 15, -8, -18, -15, -45, -11, 33, 30, 45, 43, 9, 4, 39, 96, 35, -3, -16, 16, -1, 0, -58, -22, 8, 0, 11, 64, 60, 35, -6, 0, -28, -17, 1, 29, -4, 50, 47, 67, -2, 11, -20, 59, 37, 8, 40, 59, 45, -19, -56, -21, -24, 12, 69, 52, 24, 7, 41, 29, 1, 45, -3, 8, 3, 74, 35, 32, -18, -16, -31, 62, 36, 28, 45, -36, 0, -62, -20, -2, 6, 10, 13, 29, 27, 20, 76, 36, 50, 66, 28, 19, 38, 30, 3, -6, -36, -51, -36, 62, 38, -2, 30, -9, -8, -43, -34, 8, 5, -14, 4, 2, 22, 27, 96, 57, 101, 52, 60, 15, 42, -15, -12, -18, -29, -48, -23, 40, 60, -15, 18, -22, -25, -34, -6, 33, -13, -25, -10, 38, 27, 45, 64, 64, 65, 62, 29, 16, 11, -14, -33, -28, -36, -52, -7, -2, 55, 20, -48, -55, 28, 22, 42, 35, 35, -4, -24, -27, -11, -11, 33, 37, 34, 12, 27, -25, -7, -20, -15, 2, -30, 8, -4, 28, 56, -14, -36, -23, 17, 41, 52, 39, 18, 16, -6, -16, 31, -27, -18, -16, 11, 18, 3, -17, -1, -37, 8, 12, -31, -44, 33, 57, -14, -12, -33, -32, -50, -2, 1, 10, 17, -48, -45, -43, -40, -35, -40, -22, -13, -2, -9, 1, -30, 6, -6, 22, 24, -34, -11, 12, -25, -17, -35, -71, -30, 13, 41, 36, -34, -77, -83, -79, -104, -51, -58, -25, -28, -25, -21, -74, -14, 1, -35, -11, 48, -54, -45, -34, 9, -12, -49, -33, -40, 35, 20, 28, -15, -10, -48, -90, -96, -96, -53, -61, -35, -38, -88, -116, -90, -95, -63, -72, -29, -25, -28, 5, -6, 9, 14, -15, -39, -54, -84, -37, -40, -82, -65, -135, -153, -130, -135, -160, -170, -159, -135, -87, -119, -129, -101, -75, -56, -31, -22, 6, 6, 5, -18, -18, -41, -59, -97, -119, -124, -144, -211, -166, -160, -120, -102, -101, -84, -124, -148, -105, -83, -117, -98, -55, -38, -36, -24, -12, -13, -4, 5, -10, 12, 1, -42, -64, -43, -87, -87, -126, -119, -89, -56, -11, -73, -108, -89, -60, -56, -45, -49, -32, -22, 6, 17, -9, 3, 1, -19, 20, -7, 16, -20, -15, 17, -11, -13, -4, 8, -11, -3, 23, -16, -27, 17, -19, 2, -8, 12, 0, -13, -17, -17, -7, -3, 13, 689, 6, 19, 8, 17, -41, 23, 13, 12, -8, 16, -19, -32, 8, 2, -50, 4, -28, -27, -18, -8, 11, -5, -27, -5, -19, 0, 0, -7, 1, -16, -5, -11, 11, 16, 20, 28, -9, -4, -6, -2, 41, 74, -4, 2, -13, 24, 21, -3, 47, 82, 52, 99, 25, 14, -3, -10, 18, -32, -3, 5, 29, 33, 43, 59, -6, -13, -10, -46, -47, -15, -70, -66, -41, -37, -74, -63, -48, -22, 27, -16, 18, -8, 16, 9, -16, -5, -13, -35, 56, 35, 33, 28, -20, 5, -2, 5, 0, -50, -14, -23, -22, -21, -40, -18, -12, 18, 13, -18, -92, -29, 6, -13, 14, -45, -3, -13, -21, -3, -1, 6, -9, 18, -16, 3, 27, 14, 10, 10, -4, 6, -20, 24, 11, 5, -17, -79, -20, -77, -12, 6, 8, -7, -31, -29, -51, -25, -45, -42, -29, -15, -35, 17, 25, 8, 18, 11, -13, 16, -12, 3, -17, 19, -5, -48, -27, -24, -21, -6, 3, 34, -26, -24, -63, -61, -42, -7, -21, -23, -15, 0, 3, 9, 30, 31, -4, 15, -37, 4, -49, -35, 13, -15, -71, -39, -21, -10, -2, -14, -38, -25, -51, -12, -2, -6, 4, -24, -30, -5, -27, -10, 18, 34, 10, -38, -36, -73, -39, -41, -18, -11, -54, 9, -2, 0, -12, -24, -76, -23, -6, 20, 9, 3, -9, -11, -27, -30, -32, -31, -12, 9, 8, -53, -55, -45, -36, -60, -31, -57, -64, 22, -3, 6, -43, -41, -34, -51, 5, 33, 45, -18, -12, 24, 1, 16, -36, -26, -61, -26, -38, -55, -34, -24, -16, -17, -59, -52, -104, -21, -1, -9, 12, -113, -44, -15, 6, 20, 0, -34, -17, 10, 1, 19, -1, -27, -62, -50, -41, -36, -12, 10, 16, 17, 15, -41, -97, -30, -15, -6, -52, -102, -8, 20, 17, 21, -24, 5, -2, 36, 50, 26, -16, -49, -74, -9, 32, 9, 27, 78, 132, 98, 96, 13, -45, -46, -25, -3, -50, -90, -2, 59, 51, 40, 54, 25, 38, 32, 38, 20, -4, -52, -27, 16, 94, 100, 110, 163, 162, 158, 144, 81, 15, -58, 2, -10, -37, -70, 41, 136, 139, 86, 68, 39, 24, 37, 43, 20, 13, -33, 24, 88, 111, 132, 135, 152, 185, 179, 167, 79, 22, -65, -2, -14, -28, -78, 43, 123, 144, 108, 65, 27, 35, 34, 36, 54, 52, 23, 47, 96, 111, 115, 69, 99, 127, 120, 68, 80, 32, -68, 2, 13, -29, -83, -1, 92, 138, 128, 80, 3, 12, 21, 34, 47, 47, 15, 35, 63, 56, 40, 39, 23, -20, 52, 15, -15, -28, -25, -56, -13, -13, -113, -76, 2, 24, 29, 60, -12, -2, 11, 33, 17, -18, -11, -33, -29, -5, 6, 2, 4, -14, -19, -59, -85, -48, -61, -14, -16, -37, -122, -93, -31, -29, -36, 7, -28, -22, 9, -14, 13, 3, -64, -83, -88, -40, -46, -35, -12, -2, -40, -42, -63, -69, -69, -11, -40, -8, -148, -111, -74, -52, -94, -18, -19, -1, -22, -33, -29, -22, -36, -54, -45, -37, -19, -20, -29, -25, -37, -56, -55, -89, -56, -38, -16, -57, -119, -63, -28, -70, -58, -10, -1, -36, -20, 7, 18, 20, -29, -41, -33, -15, -6, -25, -39, -54, -11, -53, -38, -71, -19, -22, 42, -23, -64, -39, -2, 13, -21, 5, 20, -17, -13, 28, 12, 51, 10, 24, 11, 45, 3, -3, -29, -16, 13, -19, -48, -70, 46, -66, -16, -5, -55, -67, -60, -16, 1, 8, 4, -2, 24, 12, 19, 40, 19, -2, -14, -2, -31, -29, 0, 6, -37, -16, -29, -46, 52, -19, 3, 36, -48, -42, -21, -20, -43, 0, -14, 24, 34, 21, -39, -38, -25, -17, -22, -40, -22, -58, -21, -26, -13, -67, 14, -22, -26, -18, 19, 25, -26, -75, -33, -11, 4, 29, 25, -16, -2, -27, -56, -63, -58, -35, -66, -50, -73, -40, 0, 11, -3, -4, -3, -33, -15, -2, 7, -4, 19, 12, 53, 32, -42, -5, -21, -19, 10, -5, 6, 10, -10, -20, -65, -12, -20, 1, 1, -8, -6, 11, 24, -6, -39, -10, 20, 1, -3, -18, -16, 4, 22, 15, 9, 4, -5, -3, 3, 30, 43, 19, 22, 56, 50, 16, 26, 37, 35, 4, 32, 21, 0, 14, 16, -12, 16, 16, 7, 12, 60, 43, 47, 27, 73, 28, 20, 18, -4, 73, 70, 48, 64, 29, 44, 50, 23, 6, 3, 2, -4, -1, -14, -12, -6, 12, 2, -20, -6, -13, 2, -1, -11, 7, 4, 18, -13, 7, 14, 15, 19, -18, -18, 4, -1, -2, 16, 2, -4, 6, -19, 80, 8, 15, 17, 1, -17, -19, -18, -19, -7, 29, 12, -36, 8, -4, -36, -7, 11, -2, -4, -37, -13, 9, -16, -11, 15, 1, -13, 0, -11, -2, 7, -11, -13, -15, -39, -41, 32, 0, -27, -76, -69, -23, -34, 35, 19, -58, -30, -30, -56, -3, 16, 51, 24, 8, 2, -13, -3, 0, 10, -20, -11, -47, -66, -23, 7, -63, -50, -67, -62, -24, -37, -18, 18, 18, -41, -96, -60, -50, -87, -70, -15, 12, -17, 3, -1, -13, -38, -28, -53, -96, -147, -83, -56, -60, -76, -24, 8, 11, 33, 59, 19, 30, 7, 13, -23, -17, 2, -33, -63, -35, -15, 1, 14, -36, -24, -43, -63, -92, -123, -85, -66, -50, -38, 12, 25, 25, 39, 23, 6, 4, 32, 57, 20, 12, 24, -28, -18, -51, -1, -9, 10, 12, -11, -65, -109, -94, -61, -74, -65, -44, -44, 11, 38, 46, 65, 32, 40, 47, 8, 25, 39, 21, 26, 0, 37, -82, -4, 16, -7, 10, -35, -74, -88, -46, 0, -7, -48, -10, -26, -41, 5, 38, 19, 35, 44, 39, 57, 17, -23, 7, -21, -4, -19, -54, -8, 20, -2, -54, -26, -59, -48, 4, 18, -36, -25, -34, -40, -39, -10, -37, -21, 22, 58, 102, 73, 8, -22, -31, -13, 44, -38, 19, 13, 9, -29, -38, -70, -26, -9, 24, 11, 20, -54, -60, -5, -17, -51, -38, -53, 7, 85, 59, 79, 20, -9, -52, -26, 35, -5, 40, -7, 11, -45, -99, -43, -28, -27, 2, 13, -2, -39, -34, -35, -16, -49, -73, -90, 18, 41, 25, 26, 7, -21, -54, -6, 4, -26, -30, -20, -30, 27, -84, -55, -30, 0, -2, 3, -11, -21, -42, -10, -36, -33, -65, -47, -21, 25, 55, 12, -19, -30, -20, 26, -2, -12, -38, -45, 8, -38, -110, -47, 3, -32, -13, 20, -11, -18, -32, -20, -66, -46, -29, -29, 16, 5, -12, -15, 14, -13, 3, 66, 8, -23, -8, -18, -23, -36, -126, -19, 21, -11, 0, 51, -9, -12, -41, -50, -63, -65, -21, 19, 28, -15, -1, -4, 10, 52, 0, 29, 4, -41, -24, -30, 40, -42, -104, -49, 19, 19, 32, 41, 9, -8, -53, -55, -38, -2, 10, 22, -12, 14, 23, 27, 19, 34, 24, 8, -52, -37, -22, -32, 15, -60, -119, -78, 26, 83, 78, 42, -10, -10, -31, -63, -31, -14, -21, 10, 2, 10, 8, 13, -6, -18, 16, -45, -76, -30, -22, 8, 0, -54, -95, -58, 54, 91, 56, 53, 39, 20, 11, -28, -42, -31, -12, 22, -3, 14, -45, 0, 4, -10, 21, -71, -118, -55, -13, -21, 14, -69, -67, -54, 75, 58, 14, 41, 7, -19, -12, -55, -51, -32, 15, 27, -7, 1, -50, -19, -50, -14, -38, -106, -132, -89, 4, 19, -14, -93, -38, -49, 48, 26, 8, -22, -10, -75, -59, -69, -77, -36, 10, 50, 38, 20, 4, -34, -53, -107, -104, -108, -87, -51, 3, 11, -23, -29, -92, -49, -16, -51, -89, -62, -48, -61, -63, -76, -57, -47, 21, 56, 67, 40, -32, -38, -98, -86, -120, -105, -63, -64, -12, -41, -23, -14, -78, -96, -45, -54, -89, -39, -35, -29, 23, -2, 1, -31, 30, 78, 75, 40, -22, -47, -120, -109, -117, -89, -70, -35, -16, -18, 24, 10, -60, -83, -51, -32, -12, -14, -6, 26, 39, 47, 17, 34, 35, 48, 27, 39, -12, -67, -163, -129, -102, -36, -31, -45, -35, -80, 1, 35, -35, -67, -72, -3, -1, 18, 22, 42, 2, -4, -16, 41, 13, 18, 1, -11, -63, -136, -127, -114, -50, -66, -53, -65, -3, -11, 0, 41, 17, -20, -23, -7, 5, 64, 54, 39, 17, -8, -38, -3, -8, -37, -50, -80, -68, -127, -154, -126, -68, -51, -60, -51, -1, -11, 20, 39, 3, -11, -15, 55, 47, 47, 41, 1, -7, -4, -16, -13, 1, -59, -85, -108, -140, -168, -151, -95, -70, -23, 13, 8, -28, 15, 1, 18, 12, 18, 40, 62, 31, 39, -16, 36, 18, 9, 12, 32, 50, 28, -49, -77, -79, -41, -42, -13, 24, 6, 29, 51, -4, 13, 14, 17, 15, -7, 18, 62, 84, 79, 77, 69, 46, 37, 22, 40, 42, 24, 22, 25, 18, -8, 10, 35, 42, 38, 51, 33, 13, -8, -14, -17, 20, 11, 19, 42, 66, 61, 82, 43, 84, 69, 33, 37, -26, 34, 58, 70, 46, 0, 28, 26, -2, 19, 23, -11, -2, -5, 17, -18, 2, -18, -7, 3, -20, 4, -19, 12, 8, 10, 5, 16, -12, 9, 6, 2, -4, -7, 9, 0, -6, 4, 5, 9, 19, 6, 9, -642, -9, 17, 7, -15, 37, -26, -7, -21, -24, -28, -7, -20, -25, -70, -43, -34, -58, -13, -41, -15, -21, -23, 12, -1, 5, -20, 0, 2, -19, -13, -8, -8, -40, -57, -107, -134, -82, -107, -24, -1, -51, -129, -43, -49, -63, -7, 9, -20, -50, -37, -28, -21, 10, -6, 1, -20, -3, 27, -2, -38, -53, -65, -103, -107, -118, -82, -27, 21, 4, 22, 31, 30, 81, 73, 39, 42, 1, -8, -3, 16, -34, -17, -6, -20, -15, 28, 49, 2, -39, 5, -15, -77, -98, -103, -30, 5, -12, 8, -4, 24, 58, 29, 51, -25, -33, -10, 0, -10, 4, 20, 18, 3, -5, 2, -50, -29, -31, -39, -38, -70, -80, -76, -66, -39, -28, -37, -22, 22, 25, 27, 0, -33, -25, -75, -62, -2, 23, 13, -17, 18, 3, -9, -45, -2, -6, -5, -31, -14, -52, -60, -81, -32, -1, -44, -11, -15, 8, 9, -45, -48, -84, -107, -43, -7, 38, 65, 0, -20, -1, 13, -19, 4, 22, -27, -12, -40, 5, -48, -44, -17, 4, -45, -26, -43, -39, -48, -75, -38, -70, -77, -23, 27, 52, 49, 48, 15, -23, 66, -26, -19, -51, -14, 41, 4, -39, -10, -22, 11, 22, -1, -25, -47, -64, -105, -102, -87, -49, -5, 17, 53, 75, -5, -39, 4, 38, 75, 2, -14, -29, 27, 67, 16, 9, 22, 50, 33, 26, 11, -36, -52, -72, -107, -65, -46, -8, 49, 50, 71, 113, -37, -3, -17, 40, 18, 62, 40, 53, 57, 56, 52, 80, 95, 39, 47, 32, 28, -14, -21, -61, -80, -33, -35, 30, 32, 37, 58, 103, 2, -10, -55, -17, 64, 121, 12, -2, 29, 61, 52, 85, 87, 58, 42, 32, 57, 15, -10, -34, -32, -21, -15, 31, 44, 31, 49, 41, 32, -24, 18, 4, 109, 49, 36, -13, 12, 53, 68, 58, 44, 63, 48, 78, 15, -31, -22, -11, 18, 25, 30, 59, 42, 32, 36, 58, -17, -22, 9, 61, 81, 22, 1, 3, 18, 21, 4, 28, 26, 44, 53, 19, -19, -36, 4, 50, 10, 36, 27, 53, 51, 41, 32, 85, 23, -7, -6, 42, 88, 36, 13, -14, -4, 0, 15, 33, 29, 18, 17, -1, -42, -36, 31, 54, 27, 34, 33, 47, 34, 26, 9, 42, -12, -37, -2, 62, 80, 64, 28, -11, -17, 50, 36, 19, 26, 23, 0, -20, -23, 11, 86, 87, 29, 13, -11, 2, -14, -35, -87, -33, 4, -34, -11, 11, -8, 20, -25, -78, 13, 7, 0, 22, 22, -47, -38, -67, -18, 64, 120, 57, -5, -54, -38, -78, -108, -105, -92, -13, 15, 0, 5, -57, -41, -29, -107, -89, -10, 14, -18, 39, 3, -49, -51, -61, -43, -34, 11, -37, -72, -101, -118, -103, -112, -99, -105, -9, -3, -31, -15, -8, -34, -18, -80, -44, 5, 4, 36, 42, 1, -56, -105, -56, -41, -18, -19, -35, -77, -86, -106, -90, -107, -55, -91, -11, -19, 27, -3, -16, -38, -55, -64, -28, 40, 35, 34, 16, -10, -85, -112, -36, 7, 11, -8, -26, -70, -64, -102, -54, -47, 0, -34, 1, 13, 11, 13, -25, -21, -3, -49, -5, 11, 31, 8, -25, -77, -124, -116, -23, 4, 39, 17, 9, -11, -31, -70, -28, 10, 37, 28, 6, -5, 0, 4, 5, 19, -26, -10, 7, 49, 15, -9, -35, -103, -80, -94, -57, 24, 51, 48, 41, -26, 8, 27, 25, 89, 55, 78, 67, 10, 37, 21, -3, 15, 7, -11, 19, 4, -14, -30, -56, -122, -100, -82, -53, 9, -8, 10, 6, -12, 73, 27, 75, 68, 75, 64, 43, 9, 2, -7, -1, -26, 43, 19, 23, -46, -53, -39, -53, -91, -106, -51, -24, -21, -11, 47, 22, 34, 59, 88, 80, 63, 57, 47, 18, 1, -13, 13, 6, -15, 36, 19, -19, -11, -18, -36, -43, -16, -60, -28, -41, -13, 19, 15, 9, 36, 28, 52, 53, 103, 72, 8, -68, -20, 0, -10, -17, 10, 35, 51, -29, -4, 16, 13, -19, -5, -3, -23, -10, -43, -54, -45, 9, 31, 24, 8, 14, 40, 9, -60, -23, -11, 18, 9, -19, 8, 25, 17, -20, -67, -8, -18, -22, -48, -35, -47, -12, -14, -2, -25, -4, 29, 42, 47, -52, -51, -3, -49, -43, 13, 20, 20, -10, -10, -13, 19, -46, -57, -61, -83, -57, -84, -69, -2, -35, -21, -66, -65, -64, -84, -70, -19, -36, -47, 8, -15, -8, -5, -15, 17, -8, 16, -3, 1, 0, -2, -8, 8, -6, -10, -16, -12, 4, -14, -17, -18, 11, 10, -13, -3, 0, 8, 4, 7, -14, 12, 11, -8, -1701, -6, -8, 0, 2, 59, 29, 28, 20, 6, 34, 68, 54, -6, -28, 34, -20, 6, 21, 14, 24, 47, 37, 11, 32, -16, 2, 14, 0, -2, -5, 12, -17, -18, 32, 20, 31, 69, 48, 9, 6, 22, 42, 57, 16, 16, 21, -21, 27, 47, -19, -26, -35, 12, -2, 6, -6, -18, -3, 10, 22, -66, 3, -14, -24, 40, 4, 35, 74, 25, 39, 11, 59, 2, -59, -43, 13, 1, 31, -13, -15, 25, -30, 3, 15, -11, 17, -3, -50, -137, -92, -83, -41, -30, -62, 18, -34, -26, 4, -25, -40, -65, -99, -71, -42, -10, -1, 10, 36, 17, 15, -20, -15, -9, 3, -41, -84, -197, -123, -145, -94, -107, -75, -75, -71, -11, -73, -74, -91, -126, -118, -104, -109, -107, -36, -22, -31, -43, -29, 5, -14, 1, 43, -17, -124, -181, -145, -161, -115, -98, -38, -43, -25, 20, -4, -37, -18, -80, -20, -2, -92, -88, -141, -94, -53, -52, -36, 7, -15, 1, 40, -44, -106, -195, -178, -134, -112, -64, 10, 33, 49, 45, 57, 35, 31, 30, 8, 21, -15, -58, -83, -108, -93, -83, -16, 7, 20, 13, 1, -71, -99, -117, -130, -82, -82, -13, 21, -5, 21, 52, 66, 39, 58, 28, 37, 9, 9, 5, -58, -55, -5, -53, -18, -42, 20, -9, -36, -48, -79, -61, -47, -22, -40, 15, 0, 3, 3, 5, 63, 42, 42, 28, -16, -14, 3, -4, 2, -36, -13, -11, 12, 28, 2, -18, 7, 27, -22, -30, 2, 19, -7, -6, 46, 1, -7, -7, 20, 58, 11, -22, -52, -28, 4, -12, -10, 17, -27, -34, 40, 18, 39, 9, -2, 28, -15, -6, 28, 29, 26, 12, 35, -13, -46, -23, 33, 7, -38, -42, -19, -43, -51, -27, 34, 5, -63, -49, 10, 5, 14, -3, -33, 7, -20, -2, 51, 94, 76, 64, 4, -46, -53, -28, 36, -21, -39, -20, -24, 1, -9, -24, 43, -3, -46, -49, 50, 15, -9, -34, -84, 38, 11, 61, 74, 93, 84, 106, 48, -39, -58, -24, 24, -9, -32, -8, -30, -34, -20, -1, 25, 11, -19, 31, 41, 2, -21, -56, -26, 49, 58, 86, 75, 54, 72, 48, 5, -31, -29, 19, 5, -39, -54, -12, 23, -15, -11, -35, 31, 6, 19, 70, 66, 12, -23, -35, -57, 5, 48, 86, 61, 64, 15, 7, 24, -2, 23, 10, 33, -43, -43, -8, 5, -20, -22, -11, 5, 34, 41, 37, 62, 16, -5, 40, -7, -16, 37, 66, 50, 8, 9, -9, 33, 36, 68, 19, 37, 35, 32, 41, 32, 13, 24, 27, -26, 25, 39, 54, 75, 38, 34, 26, -96, -72, -1, 11, 77, 36, 28, 29, 35, 3, 10, 62, 120, 104, 48, 55, 29, 0, 19, 23, -8, 43, 75, 67, 86, 43, 42, 6, -15, -70, 12, 14, 13, 17, 20, -41, -30, -42, -15, 63, 113, 114, 45, 10, 8, 6, -12, 30, 7, 37, 60, 33, 77, 27, 35, 29, -53, -113, -66, -19, 6, -7, -27, -55, -72, -67, -13, 51, 97, 41, 17, -6, -24, -1, 13, 40, 34, 56, 103, 44, 13, 67, 36, -39, -78, -173, -105, -43, -50, -52, -84, -96, -128, -89, -86, -46, -17, 11, -18, -10, 12, -18, 29, 46, 1, 29, 85, 36, 0, 58, -12, -24, -46, -131, -154, -158, -163, -109, -101, -129, -104, -141, -143, -79, -51, -43, -35, -5, 14, 0, -28, 43, -7, 28, 47, 61, 1, 24, -7, -34, -48, -90, -188, -227, -197, -120, -103, -105, -86, -122, -91, -101, -74, -65, -49, -26, -30, -21, -36, 4, -24, 24, 67, 42, -19, 18, -19, 23, -19, -81, -114, -90, -111, -67, -74, -49, -33, -82, -54, -40, -64, -28, -68, -51, -33, -31, -23, -28, -19, 2, 69, -59, 53, 18, -19, -12, -10, -59, -78, -14, -44, 9, 2, 23, -8, -50, -17, -30, -2, 3, 3, -15, -2, 15, -3, -22, 13, 13, 63, -4, -7, -15, 13, 14, -5, -40, -10, 10, 50, 68, 58, 60, 30, 24, 23, 52, 26, 71, 36, 35, 12, 84, 72, 54, 55, 36, 41, 5, -4, -6, 2, 9, 19, -27, -2, 72, 76, 124, 82, 56, 49, 27, 31, 71, 21, 13, 50, 79, 31, 30, 27, 60, 31, 15, 49, 16, 3, 2, -6, -17, -5, -16, 18, 58, 51, 58, 70, 67, 66, 44, 33, 44, -32, -7, 63, 31, 31, 39, 23, 34, 37, 28, 13, -9, -2, -18, -3, -17, -2, 8, 12, -11, 16, 7, 0, -19, -20, 14, -3, -15, -23, 21, 24, 4, -2, -6, -7, -1, 9, 15, -20, -10, -9, -12, 14, -1873, -13, 9, -15, -10, 41, -39, -45, -21, -28, 1, 42, 31, 8, -1, 39, 33, 33, 51, -4, 10, 10, 6, 3, 2, -2, 9, -15, -2, 2, -17, -12, -9, -37, -22, -13, 21, 39, 21, 4, 41, 71, 27, 37, -3, 2, 14, 18, 38, -33, -46, -64, -43, -22, 18, -2, -10, 8, 25, 2, 44, 13, -20, -43, -11, -21, -22, -40, 16, -5, 3, 8, 82, 42, 61, 90, 73, 20, 32, 8, 13, -13, -4, -9, 6, 13, 3, 22, 13, -28, -46, -25, -61, -79, -63, -7, -24, -1, -23, -33, -11, 12, 13, -1, 2, 40, 40, 30, 83, 47, 47, 5, 11, -12, 36, 5, 38, -5, -18, -35, -26, -44, -21, -7, -16, 11, -28, -39, -67, -48, -34, -16, -46, -18, 20, 47, 67, 34, 43, -12, 0, -10, -12, 9, 42, 4, -23, -23, 2, -2, -18, -2, -14, -10, -43, -34, -67, -55, -56, -86, -68, -50, -50, -32, 13, 2, 6, -3, 3, -23, -13, 54, 24, -42, -36, -15, 10, 3, 2, -17, -13, -41, -21, -52, -34, -67, -33, -54, -52, -40, -16, -24, -22, 53, 50, 11, -12, -2, 27, 62, -3, -59, -69, -21, 5, 29, -4, -42, 4, -2, 0, 2, -36, 1, 7, 3, 18, -17, 12, 25, 11, 34, -24, -15, 14, 34, 14, 131, 41, -65, -43, 34, 35, 57, -3, 14, 16, -3, 5, -22, -23, 11, 25, 43, 26, 9, 28, 5, 15, 54, -6, -28, -18, 30, 74, 68, -9, -31, -31, -12, 41, 56, 15, 10, 22, -4, -8, 1, -3, 2, 29, 10, 34, 46, 35, 60, 13, 63, 15, 33, 20, 13, 86, 3, 26, -21, -39, -39, 14, 36, 10, -1, -6, -9, -10, 15, 19, -15, -7, 27, 22, 58, 81, 48, 44, 55, 19, 28, -19, 50, 69, 41, 47, 16, -28, 1, -10, 50, 5, -19, -46, -43, 20, 25, 32, 17, 39, 46, 68, 74, 82, 67, 41, 4, 34, 33, 0, 31, 64, 26, 53, 9, -22, 14, -23, 3, 6, 0, -2, 15, 34, 61, 41, 34, 59, 48, 69, 64, 78, 47, 9, -67, -18, 21, -9, 1, 39, 15, 7, -54, -70, -32, -18, -50, -7, 5, -8, 28, 67, 56, 63, 8, 30, 34, 9, 12, -18, -67, -88, -62, -1, 3, -14, 8, 87, 21, -53, -88, -85, -43, -51, -27, 28, 25, -8, -30, 38, 33, 7, -15, -43, -98, -139, -151, -158, -195, -172, -84, 4, 1, -20, -10, 83, -6, -106, -101, -54, -89, -32, -38, -21, 1, 6, -3, 30, -55, -124, -128, -154, -192, -221, -210, -145, -132, -122, -81, -45, 3, 23, -8, 53, 54, 3, 11, 21, -38, -17, -22, -19, -15, 10, -15, -73, -163, -228, -188, -158, -155, -124, -94, -68, -63, -57, -14, -8, -22, 19, 29, 86, 115, 52, 62, 47, 18, -1, -42, -23, -9, -17, -75, -106, -119, -130, -70, -3, -19, -4, -17, -3, -43, -27, 48, 32, 8, 15, 31, 94, 86, 16, 70, 59, 9, 25, 5, 16, 33, -7, -46, -14, -40, 24, 54, 50, 57, 45, 56, 23, 1, 26, 51, 53, 47, -2, 25, 51, 29, 10, 23, 59, 22, 63, 20, 21, 30, 37, 48, 36, 73, 77, 92, 78, 36, 37, 20, -45, -26, 8, 55, 24, 26, -14, -32, 1, -19, -19, 11, -10, -34, 34, 18, 8, 7, 15, 19, 77, 48, 31, 49, 36, 34, -12, -34, -21, -26, -17, 40, 29, 71, -3, -38, 4, -44, -5, -14, 1, -12, -8, 14, -6, -15, 12, -1, 11, -12, -10, -4, 2, -15, -40, -29, -6, 34, -2, 29, 61, 36, -3, -31, -23, -77, -28, -9, 2, -23, 7, 7, -17, -51, -4, -15, -74, -75, -67, -67, -42, -44, -70, 14, -4, 24, 8, 38, 20, 1, 1, -23, -30, -7, -11, -61, -19, 7, 18, 43, 54, -27, -19, -29, -86, -89, -66, -56, -50, -101, -30, -10, 2, 3, 22, 41, 58, 21, 7, 8, -37, -50, -32, -78, -78, -35, 39, 70, 80, 70, 47, 54, 12, 44, 44, 9, -17, -7, 38, 5, -62, -25, 22, 51, 42, 16, 12, 1, -17, 21, -5, -19, -50, -33, -3, 25, 49, 66, 56, 24, -17, 2, -12, -5, 8, -1, -47, -36, -37, -10, -13, -21, -10, 16, 5, 6, -11, 18, 16, -21, -2, -32, -45, -61, -76, -48, 19, 6, -12, -70, -39, -50, -46, -36, -28, -10, 4, 5, -10, -14, 5, -14, -20, 4, -13, -11, -10, 7, 3, -2, 6, -4, -3, -8, -3, -11, -11, 1, -11, -11, -6, 11, -7, 4, -9, 7, 5, 13, 4, -13, 7, -1174, 15, -15, 13, 19, 38, 26, -2, 38, 35, 29, 41, 16, 8, 14, 81, 26, 46, 50, 66, 34, 51, 15, -7, 20, 5, -16, 13, -18, 5, 6, 2, -24, -12, 9, 21, 71, 93, 11, -18, -4, -9, 33, -20, -36, -32, 1, -13, 59, 32, -5, 12, -52, -22, 17, -11, -4, -16, 38, 52, 5, -20, -21, 16, 41, 38, -3, 0, -18, -27, -26, -48, -48, -72, -123, -89, -31, -35, -8, 23, 25, -11, -45, 20, 10, 12, 28, 64, 95, 45, 25, 54, 1, 51, 29, 8, -16, -38, -19, -68, -67, -64, -71, -21, -34, -1, 25, 22, -14, -83, -5, 4, -15, -13, -18, -15, -2, 46, 21, -3, 17, 3, 17, 29, 5, 15, -24, -8, -23, -17, -5, 16, 9, 29, 59, 55, -22, -86, -19, -12, -20, 3, -39, 6, 64, 43, 26, 1, 34, 29, 54, 21, -28, -15, 8, -5, -15, -25, 8, 34, 51, 61, 27, 52, 19, 12, 34, -20, -16, -8, -32, 10, 55, 47, 19, -1, -3, 38, 40, -3, 34, 36, 7, -10, -12, -23, 27, 25, 24, 2, 6, 41, 33, 16, 10, -3, -17, -11, 65, 48, 39, 9, -8, -5, -13, -30, 4, 19, 34, 32, 37, -11, 0, -4, -4, -6, 29, 29, 30, -13, 23, -12, -36, -33, 13, 32, 42, 33, -11, 4, -13, -30, -26, -34, 16, 12, 22, 45, 7, 19, 7, -3, 29, 20, 19, 8, 6, -45, -9, -38, -31, 6, 18, 38, 43, 41, -7, 15, -6, -48, -28, -9, -15, 9, -12, 49, 15, 13, 14, 9, 14, -16, -27, -22, -33, -26, -48, -53, -19, -18, 12, 60, 88, 81, 5, -26, -42, -33, -29, -8, -7, -4, -9, 34, 68, 43, 30, -1, 7, -18, -59, -97, -103, -115, -85, -65, -26, -17, -10, 67, 76, 14, -2, -19, -32, -19, -29, -30, -22, 24, 11, 4, 43, 36, 11, -60, -78, -103, -140, -103, -86, -105, -70, -63, -11, -32, 0, 45, 76, 17, -42, -64, -61, -30, -12, -22, -15, 27, -16, -7, 0, 14, -56, -120, -189, -155, -130, -114, -73, -112, -83, -31, 5, -49, -26, 58, 107, 43, -56, -38, -53, -40, -47, 17, -2, 5, -17, -12, -53, -64, -126, -186, -174, -143, -128, -89, -69, -58, -74, -25, 74, -10, -6, 34, 90, 50, -24, -72, -81, -61, -48, -31, -19, 12, -15, -43, -45, -112, -178, -169, -93, -60, -54, -48, -4, -28, -10, -34, 83, 26, -17, 34, 27, 41, -36, -94, -83, -31, -28, -9, 0, -10, -9, -53, -54, -144, -107, -53, -17, -7, 36, 14, 8, 39, 16, -55, 65, 36, 21, 18, 0, -8, -94, -77, -19, 12, -5, 3, -17, 2, -19, -9, -62, -59, -5, 57, 68, 57, 50, 52, 44, 71, -17, -8, 44, 16, 29, 43, -13, -43, -53, -78, -23, 10, 13, 5, 4, -11, -30, -35, 1, 47, 55, 94, 115, 76, 53, 12, 31, 53, -31, -15, 0, -2, 12, -1, 29, -28, -66, -15, -1, 7, -7, -19, -35, -3, -59, 10, 45, 52, 82, 45, 46, 30, 6, 6, 2, 28, 6, 3, 15, 36, 10, 19, 5, -80, -95, 9, 26, 29, 26, -2, -27, -30, -23, 6, 74, 59, 41, 36, 48, -12, 31, -21, -32, -34, 13, -11, 3, 47, -16, -7, -27, -93, -51, -35, 8, 18, 16, -22, -31, -29, -2, -20, 32, 25, 21, 9, 10, 19, -9, -21, 25, -48, 25, 64, 3, 33, 8, 10, -30, -64, -49, 6, 6, 10, -7, -16, -27, 4, 9, -12, 34, 27, 34, 37, 33, 15, 1, -17, 30, -11, -2, 23, 8, -11, 10, -27, -38, -18, -21, 18, 25, -1, -4, 27, -15, -39, -23, -40, -15, 7, 23, 11, 12, 26, 21, 4, 12, 27, 30, 3, 42, 14, -20, -12, 9, -26, -62, -25, -28, -30, -17, -54, -47, -67, -83, -71, -38, -18, -52, -53, -39, -13, 14, 12, 49, 10, -33, -13, 38, 20, 15, -6, -11, 2, -47, -24, -66, -102, -76, -53, -84, -63, -73, -79, -115, -106, -68, -83, -92, -37, -60, -54, 11, 8, -23, 7, 6, 8, 11, -18, -5, 39, 43, 5, -17, -16, -73, -96, -58, -57, -60, -66, -42, -73, -44, -39, -26, 1, 34, -1, -12, -16, -2, 0, 3, 14, 18, 11, -8, -5, -10, -30, -46, -41, -40, -13, -34, 2, 9, 3, -5, -58, -68, -20, -48, -3, -23, -28, 3, -13, 16, 9, 2, -7, -19, 18, 19, -9, -9, -9, -11, -2, -1, 8, -18, -14, -17, -1, 3, -20, 12, 6, 10, 1, 6, 17, -4, 7, 9, -16, 11, 12, 20, -532, 10, -7, 15, -3, 18, 29, 55, 45, 61, 51, 49, -2, -13, -31, 31, -12, -16, 13, 3, -12, 4, -29, 19, 32, 16, -10, 16, 18, 9, 20, 20, 6, -6, -2, 38, 28, 2, 0, -26, -2, 29, 25, 3, -29, -51, 7, 40, 47, 22, 25, -28, -18, -5, -4, -8, -18, -1, 5, 27, -69, -63, -11, 33, 38, -14, 43, 21, 24, 35, 34, 3, 13, 2, -4, 1, 27, 14, 10, 22, 27, 22, -23, 8, 20, -4, 8, 75, 1, -23, 10, 22, -11, -21, -19, 15, 6, -26, -20, -32, -27, -3, 0, 23, -2, 7, 22, 25, -28, -87, -15, -20, 9, 10, -54, -59, -29, -39, -51, -23, -70, -59, -62, -78, -62, -30, -19, -61, -16, -10, -33, -33, -21, 19, -11, -52, -56, -68, -41, 10, -19, -21, -36, -25, -10, -56, -71, -82, -52, -76, -78, -72, -45, -36, -47, -72, -59, -29, -31, -47, -32, -47, -92, -58, 0, 14, 34, 12, 9, -11, -24, -19, 43, -1, -75, -59, -69, -50, -61, -22, -20, -60, -28, -31, -62, -69, -46, -41, 15, -65, -59, -16, -7, 28, 54, -2, -13, 1, 48, 36, 33, -39, -97, -43, -25, -15, -50, -23, -3, -3, 33, -12, -52, -70, -69, -42, -9, 1, 8, 33, 62, 43, 28, -54, 20, -10, 57, 20, -59, -40, -14, -27, -6, 46, 23, 54, 91, 79, 76, 6, -61, -17, -50, -61, -14, 39, 17, 68, 97, 62, -10, 30, -9, 48, 53, 52, 2, -14, -16, 42, 56, 115, 122, 103, 108, 64, 68, 15, -48, -79, -96, -44, -9, 16, 22, 42, 83, 55, -18, -16, 6, -50, 69, 106, -4, -17, -2, 83, 86, 110, 124, 81, 78, 87, 49, 0, -57, -54, -25, -21, 32, 22, 28, 22, 41, -28, 26, -50, 19, -42, 109, 50, 0, -23, 56, 92, 111, 84, 53, 61, 63, 120, 10, -68, -65, -39, -42, -1, 3, 68, 38, 32, 18, -11, -24, -57, 25, 60, 89, 1, -2, 4, 114, 63, 92, 94, 47, 36, 33, 63, -9, -71, -103, -44, -26, -1, 3, 25, 11, 11, 14, 30, -1, -36, -1, 48, 53, 45, 27, 37, 101, 56, 52, 38, -5, 34, 53, 21, -39, -99, -46, -29, 0, -5, 19, -4, 28, 40, 56, 15, 66, -1, -12, 60, 51, 32, 31, 54, 41, 55, 16, 13, 4, 23, 57, 32, -68, -101, -56, -9, 7, 4, 9, -12, 22, 24, 21, -17, 106, 24, -8, 35, -42, -24, -14, 27, 25, 31, 17, 12, 14, -15, 41, -31, -78, -93, -12, 23, 23, -4, 18, 30, -21, 6, -16, -32, 76, 62, 18, 1, -79, -47, -45, 0, 11, 21, 33, 31, -5, -30, -34, -84, -120, -63, 9, 14, 22, 6, 3, -6, 3, 4, -13, -1, 84, 30, 12, -15, -63, -14, -85, -32, 19, 17, 9, 30, 0, -20, -90, -97, -74, 7, 5, 17, 4, -5, -22, -13, 5, 6, -50, -3, 5, 69, 22, -23, -53, -38, -46, -36, -9, 18, 30, 16, 15, -28, -78, -66, -28, -13, 20, -15, -9, -22, -13, -13, -26, 20, 22, 40, 13, 63, -9, -48, 0, 32, -29, -23, -5, 13, 12, -10, 4, -58, -55, -57, -1, -5, 2, 18, 11, -5, -24, -11, 25, 42, 19, 39, 59, 54, -42, -54, 42, 33, 27, -38, -45, -10, 10, -6, -6, -1, -25, -37, -29, 22, -16, -24, -22, -18, -16, 34, 75, 20, 34, 55, 34, 17, -14, -29, -46, -5, -66, -43, -42, -25, -18, -13, -18, 7, -23, -34, -45, -43, -17, 4, -25, 46, 65, 91, 64, 63, 32, 11, 15, -18, 18, -9, -66, 57, 0, -39, -82, -103, -68, -36, -2, -20, -47, -67, -60, -22, 8, 9, 9, 53, 91, 56, 86, 44, 51, -74, -4, 5, -13, -17, -27, 43, 10, -11, -19, -50, -76, -95, -29, -50, -23, -56, -29, 0, 9, 4, 5, 35, 39, 61, 96, 57, 0, -55, -16, -11, -15, -19, 11, 67, -6, -10, 56, -11, -34, -36, 5, 13, -24, -25, -44, -72, 1, 32, 46, 32, -18, 15, 32, 27, -32, -29, 5, 13, -2, -6, 9, 22, 29, 21, -12, 46, 16, 11, -2, -7, -2, -22, -15, 4, 63, 76, 95, 96, 51, 9, 26, -7, -17, -8, 10, 7, -20, 14, 13, 4, 16, -43, -50, -58, -64, -43, -52, -17, -32, -32, -34, -3, -24, -6, 24, 32, 8, 7, -25, -12, 4, -5, 4, -14, -1, -1, 16, 2, 18, 12, 15, 17, -11, 17, -14, 20, -3, -14, -12, 9, -6, -12, 15, 12, -12, -4, 1, 4, -14, 14, 20, 19, -14, -508, -11, -6, 14, -16, 45, -4, 13, 33, 26, 38, 65, 29, -4, 2, 87, -8, 21, 40, 28, 66, 27, 38, 30, -6, 10, -7, 7, -5, -1, -15, 5, -33, -8, -2, -21, 14, 46, 16, -43, -38, -21, -6, 10, -1, -22, -4, -3, 4, 17, -28, -49, -71, -19, -6, 2, -17, -2, 25, -26, 37, -28, -14, -25, -58, 1, -6, -16, -28, -19, 7, -22, 6, -2, -37, -6, 4, 4, -27, 9, 15, 56, -36, -19, 19, -5, 43, 20, -26, -93, -73, -95, -75, -64, -99, -66, -74, -46, -35, -47, -37, -18, -19, -28, -48, -73, 5, -13, -2, -20, -23, 4, 9, -17, 7, -22, -61, -149, -138, -117, -79, -49, -91, -71, -47, -53, -53, -79, -80, -72, -54, -38, -57, -45, -17, -16, -56, -89, -53, -4, 15, 8, 51, 40, -27, -128, -154, -96, -29, -30, -23, -13, -11, 0, -12, -39, -10, -26, -14, -2, -27, -42, -44, -34, -7, -54, -26, 10, -8, -19, 39, 24, 8, -53, -100, -77, -21, -1, -3, 30, 19, 42, 79, 60, 44, 58, 49, -15, -30, -39, -72, -59, -46, -61, -3, 5, -2, 17, 41, 18, 9, -57, -60, -64, -8, 13, 22, 29, 10, 44, 80, 98, 110, 86, 18, -51, -61, -85, -103, -104, -71, -17, 1, 3, -14, 10, 23, 5, -35, -40, -16, -22, -12, -12, 3, -3, -9, 27, 91, 113, 99, 43, 11, -66, -68, -60, -41, -122, -102, -51, 31, 25, 5, 11, 62, 57, 6, 15, 5, 23, -21, -65, -17, -32, 13, 16, 54, 83, 48, -29, -47, -99, -89, -43, -59, -76, -96, -79, 15, 12, 52, -19, 47, 103, 37, -16, 10, 32, -11, -33, 3, 9, 0, 30, 79, 60, 22, -18, -57, -94, -88, -79, -61, -42, -75, -85, 1, 6, -18, -19, -31, 22, -14, -26, 25, 17, -9, 4, 8, -17, 25, 45, 51, 17, -25, -39, -79, -72, -75, -63, -19, -27, -40, -48, 15, -24, -9, -25, -69, 23, -35, 34, 57, 16, 9, 33, 1, -11, -13, 25, 38, 6, -30, -56, -61, -87, -81, -52, -21, -44, -40, 28, 71, -31, 1, 20, 0, 16, 26, 98, 87, 51, 35, 25, 9, -5, 10, 14, -1, -57, -72, -54, -36, -47, -41, -62, -4, 17, 6, 68, 72, 24, 19, -26, -25, 26, 46, 72, 53, 26, -42, -6, 13, 19, 38, 7, 1, -89, -107, -90, -60, -47, -26, -7, -7, 29, 64, 62, 91, 40, 20, 45, 2, 21, 47, 101, 55, -17, -10, -22, 22, 33, 42, 19, -7, -96, -107, -70, -36, 1, 54, 59, 17, 40, 75, 57, 35, 72, 32, 1, -91, -73, -5, 54, 49, 34, 17, -8, 17, 44, 54, 40, 32, -14, -60, -37, -29, -20, 10, 41, -14, 29, 87, 34, 72, 55, 39, -9, -14, -68, 7, 16, -19, 28, -33, -1, -3, 6, 13, 36, 41, 39, -14, 10, -28, 5, -6, 25, 43, 56, 90, -15, 40, 29, 29, 27, -44, -83, -35, -15, 26, -9, -42, -23, -29, -26, -27, -18, 26, -8, -2, 6, -10, 46, 48, 65, 39, 58, 83, 42, 42, 70, 15, -33, -85, -132, -54, -17, -10, -42, -42, -49, -64, -50, -87, -46, -48, -37, 7, 30, 41, 43, 64, 49, 53, 16, 40, 39, 37, 78, -11, -11, -66, -72, -87, -140, -93, -52, -70, -65, -47, -59, -44, -46, -38, -16, 11, 67, 44, 36, 9, 77, 32, 24, 66, 44, -2, 28, 8, -26, -42, -78, -147, -184, -143, -101, -115, -89, -78, -87, -63, -32, -35, 1, 31, 21, 33, -19, 4, 28, 57, 25, 30, -21, -6, -18, 5, 19, 8, -66, -80, -135, -132, -129, -104, -137, -101, -90, -80, -28, 2, 2, -28, -32, 14, -6, 7, -1, -8, -22, 26, -61, 8, 10, 5, 0, 30, -40, -59, -61, -68, -38, -35, -32, -60, -18, 5, 13, 58, 66, 11, 2, 7, -6, -34, -30, -66, -23, 5, 15, -2, 7, 6, 16, -3, -1, -13, 12, 14, 11, 27, 60, 7, -8, 42, 50, 75, 62, 55, 30, 23, 83, 28, 23, 35, 45, 21, 33, -23, -20, 18, 10, -1, 3, -4, 44, 44, 43, 98, 89, 61, 56, 54, 108, 99, 54, 77, 73, 60, 41, 67, 68, 89, 42, 27, 29, 16, -2, 0, 19, -19, -20, 8, 22, 41, 62, 56, 68, 100, 87, 70, 79, -2, 57, 26, 40, 40, 31, 29, 33, 64, 29, 18, -20, 7, 4, -13, -10, -6, 17, -9, 7, -7, -11, 20, 16, -15, -11, 3, -19, -21, 25, 26, -4, -2, 5, -6, 15, 4, 18, 15, 1, -3, -4, 10, -1636, -2, 0, -20, 17, 3, -36, -50, -17, -17, -32, -44, -31, -42, -82, -38, -28, -26, -30, -20, -33, -29, -24, -4, 12, -17, -19, -3, 6, 13, 7, 20, 2, -30, -61, -73, -61, -132, -127, -123, -141, -118, -134, -148, -193, -88, -115, -92, -79, -35, -41, -45, -51, -4, 14, 3, 7, 15, 18, 29, -24, -50, -56, -59, -81, -134, -185, -217, -250, -222, -196, -207, -175, -144, -122, -127, -104, -64, -81, -86, -25, -16, -17, 15, -10, 2, 13, 37, -40, -76, -18, -26, -44, -50, -60, -75, -102, -117, -130, -143, -140, -104, -75, -97, -94, -47, -29, 1, -56, -59, -16, 13, -4, 13, 49, -7, -40, -88, 7, -16, 2, 26, 1, -5, -9, -25, -74, -44, -24, -65, -37, -65, -68, -47, 18, 49, -11, -54, -4, 16, -1, -22, -9, -31, -6, -20, -34, 54, 89, 59, 60, 50, 8, -23, -35, -29, -45, -27, 8, 6, 24, -15, 6, 98, 92, 26, -17, -20, 5, -13, 24, 21, 58, 27, 11, 61, 83, 78, 86, 28, 5, -11, -6, -46, 7, -25, -3, 18, 7, -1, -11, 40, 86, 21, -4, 3, -5, 0, 78, -12, 26, 37, 18, 50, 74, 52, 68, 29, 24, 1, 3, -28, 7, 9, 6, 28, 49, 33, 17, 0, 38, -13, 6, -22, 21, 27, 71, 51, 32, 58, 43, 36, 37, 66, 38, 4, 7, 26, -8, -18, 13, 7, 22, 48, 52, 37, 12, -4, 42, -1, -15, -50, 19, 34, 1, 94, 32, 59, 55, 74, 28, 43, 13, -27, -8, 13, 51, 35, 45, 29, 52, 56, 55, -3, 7, 38, 44, 51, -22, 3, -20, 11, -1, 69, 29, 35, 52, 42, 32, -9, -11, -24, 12, 31, 74, 54, 52, 43, 83, 44, 19, 16, 23, -1, 15, 3, -19, -25, -18, 17, 47, 87, 29, 47, 57, 13, -9, -35, -28, -17, 42, 46, 69, 65, 67, 80, 65, 48, -24, 20, 8, 11, -6, 39, -27, -39, 0, 41, 37, 82, 33, 7, -1, -27, -32, -64, -51, -50, 6, 52, 79, 83, 61, 25, 11, -1, 14, 16, 1, -26, 8, 40, -2, -54, 18, 59, 92, 53, -17, -33, -16, -44, -61, -60, -52, -43, 23, 15, 30, 27, -21, -43, -51, -9, -17, 13, -1, -39, 1, 43, -43, -60, 4, 41, 42, 18, 1, -21, -9, -15, -47, -24, -57, -44, 4, 15, 22, 41, -35, -36, -15, -28, -14, -28, -19, -35, -67, -46, -22, -12, 8, 45, -54, -1, -36, -18, 22, -5, -21, -34, -35, -85, -16, -14, 2, -5, 10, -33, -19, -10, -36, -46, -47, -23, -70, -107, -24, -22, 15, -33, -80, -40, -136, -64, -8, -11, -34, -24, -114, -97, -42, 11, 9, -11, -22, -3, 12, -30, -46, -32, -50, -32, -45, -93, -18, 8, 6, -13, -46, -68, -125, -107, -58, -55, -71, -74, -123, -86, -40, 8, 34, 5, -6, 6, -23, -57, -53, -36, -27, -30, -92, -90, -38, -17, 12, -7, -45, -117, -138, -92, -53, -49, -49, -97, -138, -104, -57, 13, 33, 18, 21, 4, -10, -37, -77, -48, -76, -72, -88, -18, -33, -53, 14, -21, -35, -111, -123, -71, -40, -30, -37, -34, -79, -41, -51, -4, 26, 19, 18, 13, -25, -67, -98, -93, -80, -85, -85, -80, -10, 40, -24, 15, -2, -68, -49, -44, -5, -2, 23, -25, -51, -12, -24, -12, 15, 35, 32, 15, -18, -95, -102, -87, -90, -124, -92, -96, 1, -4, -18, 4, -10, -4, -12, -33, -19, 15, 7, 0, -4, -24, -11, 23, 12, 17, -26, -17, -65, -119, -130, -66, -58, -71, -49, -56, -22, 5, -18, 19, -2, -4, 66, 31, 23, 39, 34, 32, 29, -15, 24, 51, 20, 3, -39, -59, -85, -95, -40, -25, -4, -8, -18, -14, 42, -19, 17, -26, -81, -48, -36, 19, 6, 29, 16, 16, 0, 9, 25, 13, -2, 8, -65, -71, -42, -46, -9, -5, 33, 33, 19, -44, 7, -21, 11, -15, -10, 18, 25, -1, 9, 17, -51, -43, -41, 15, -2, 4, -26, -17, -95, -82, -35, -9, -9, 15, 28, -11, 5, -7, 12, 16, 9, 5, -9, 22, 80, 35, 34, 56, 36, 28, 35, 47, 42, 153, 119, 88, 97, 109, 113, 131, 106, 78, 50, 0, 6, -9, 26, -1, 12, -18, -11, 5, 19, 21, 55, 25, 65, 53, 90, 29, 2, 40, 23, -7, 16, 28, 75, 64, 31, 54, 21, 20, -18, 9, -4, -3, -7, 17, 18, -13, -2, -8, -9, 9, 17, 7, 19, 17, -14, 5, 4, 2, 12, 1, -19, -6, -1, -2, 4, 17, -17, -6, -1, 10, -11, 85, -5, 1, -16, -9, 27, 10, -11, -24, -15, -18, 0, -4, -27, -29, 20, -1, -2, 11, 5, 27, 11, -4, -2, 20, 12, 6, 12, 12, 2, 5, 17, -31, -41, -34, -37, -64, 10, 16, -5, -47, -31, -37, 9, 8, 7, 43, -16, -28, -24, -61, -49, -62, 11, 10, -19, 0, -19, -36, -7, 42, -9, -55, -77, -55, -14, 7, 25, 25, 15, -4, 35, 65, 65, 102, 71, 80, 98, 60, -18, 39, -30, 1, 4, 15, 1, -3, -50, -26, -30, -51, -62, -63, -29, -38, -46, -24, -34, 4, 30, 14, 39, 56, 13, 21, 15, 47, 39, 51, 58, 39, -9, 15, -10, 55, -13, -34, 1, -21, -36, 17, -9, 5, -34, -25, -21, -51, 5, 14, 26, 39, 17, 23, 4, 13, -5, 34, 53, 68, -10, -6, -16, 16, 20, -30, 9, -10, 18, 33, 18, -4, -16, -38, -28, -23, -23, 4, 12, 8, 52, 7, 2, 10, -12, -30, -39, 8, -12, 14, 1, -65, 15, -50, 23, 5, 13, 33, 31, 34, 1, -37, -5, 20, 18, 25, 24, 15, 24, 37, 44, -5, -52, -43, 6, -14, 7, 17, -19, -64, -22, -16, 34, 39, 53, 43, 4, -11, -13, -44, -42, 9, 46, 39, 17, 37, 32, 54, 47, 1, -26, -56, -4, -44, -24, -15, -11, -25, -13, 23, 32, 29, 32, 23, -28, -18, -30, -94, -62, -17, 79, 83, 20, 20, 12, 8, 4, -1, 25, -22, -10, -29, 16, -18, -11, -19, -64, 32, 50, 24, -9, 11, -33, -51, -73, -122, -97, 37, 118, 87, 52, 8, -12, 16, -12, 23, 26, 1, 62, 52, 20, 19, -27, -41, -41, 45, 51, -32, -25, -28, -33, -75, -94, -95, -56, 90, 137, 82, 12, -28, -10, -31, 7, 8, -23, 13, 60, 5, 49, 9, -20, -14, -11, 39, 22, -52, -18, -31, -51, -73, -107, -67, 19, 112, 128, 27, -8, 20, 30, -4, -26, -34, -30, 7, 51, 33, 34, -14, -23, 12, 1, 24, -20, -22, -37, -10, -43, -52, -86, 2, 50, 102, 66, 25, -13, -12, -8, 4, -51, 0, -75, -44, -12, 30, 40, 22, 12, 21, -13, -8, -41, -50, -20, -50, -27, -28, -19, 21, 85, 89, 42, 3, -28, -42, -20, -30, -68, -23, -46, -86, -27, 52, 19, 4, 37, 38, 20, -23, -38, -66, -41, -25, -20, -16, -18, 42, 59, 60, 19, -39, -13, -54, -37, -29, -44, -18, -32, -79, 5, 23, -7, -14, 44, 68, 71, 16, -24, -43, -8, -11, -24, 1, -4, 15, 95, 98, 42, 6, -38, -33, -24, -30, -10, -6, 31, 2, 43, -2, 12, -5, 30, 92, 88, 76, 36, 25, 5, -8, -38, -13, 12, 11, 65, 113, 45, 14, 11, -1, -6, -11, -8, -18, 7, 18, 61, 44, -13, -10, 16, 46, 68, 65, 57, 25, 0, 2, 6, 7, -20, 40, 68, 67, 58, 1, -36, 9, 4, 15, 19, 6, -46, -10, 43, -3, -9, 42, 8, 55, 84, 63, 61, 75, 64, 28, 34, 6, 20, 34, 50, 31, 37, 16, -18, -32, -3, 0, 11, 1, -22, 20, 23, 45, 31, 9, 41, 15, -12, 21, 80, 78, 22, 34, 39, 39, 34, 26, 14, 3, 25, 12, -13, -7, 1, -16, 4, -15, -55, 7, 42, -19, 19, -45, 18, -8, 12, 13, 83, 74, 24, 12, 24, -1, 18, 35, 10, 12, -8, -2, -20, -24, -24, 13, 4, -26, -29, 0, 25, -43, 80, 5, 40, 30, 77, 49, 46, 59, 54, 25, 20, 30, 39, 27, 8, -13, -13, -6, -3, 4, 16, 9, 30, 8, -4, -18, 26, -15, 26, -2, 11, 65, 60, 35, 30, 11, 15, 52, 0, 2, -6, 23, -18, -3, -36, 19, 0, -17, 7, -5, 32, 34, 23, 8, 27, 11, -8, 11, 25, 32, 8, 30, -32, -67, -23, -4, 10, 19, 16, 39, 30, 16, 17, 41, 39, 59, 39, 46, 14, -11, 14, 42, 66, 31, 6, 10, -18, -4, -19, -15, -20, -1, 0, 53, 26, 50, 8, 21, 6, 12, -22, 1, -4, -4, -14, -15, -21, -36, 7, 24, 40, 15, -13, 12, -8, -6, 35, 20, 23, -13, -15, -2, 3, 47, 29, 12, -15, -39, 13, -43, -21, -67, -64, -60, -50, -56, -5, 32, -28, 5, 12, -9, -6, 3, -10, -12, 3, 7, 41, 37, 12, 15, -23, -17, -7, -6, -22, -51, -24, -22, -14, -6, 4, 34, 11, -3, 6, -1, 4, -16, -9, 4, 10, -9, -7, 18, -2, 7, 20, 15, -2, 10, 9, -17, -10, 0, 7, 9, -18, -4, -11, -10, 11, -1, 20, 6, 0, 12, 247, -4, -13, -19, 3, -55, -43, -16, -29, -27, -27, -70, -50, -18, 7, -40, 11, -10, -27, 0, -29, -50, -24, -21, -17, -13, 13, -5, -14, 4, -2, 0, -5, -33, -67, -39, -43, -92, -72, -102, -99, -106, -75, -85, -18, -49, -46, -1, 20, 47, 32, 49, 82, 18, -9, -15, -3, -1, -9, 2, -13, 6, -39, -28, -4, -17, -12, 5, -51, -53, -32, -27, -77, -71, -91, -110, -114, -67, -35, -63, -34, -56, 10, -9, 14, 2, -18, 18, 51, 88, 86, 77, 73, 73, 52, -1, 25, 30, 14, 35, 33, -2, 8, 24, 11, 18, -6, -92, -60, -89, -19, -3, -2, 11, -25, 15, 28, 93, 113, 93, 75, 67, 12, -5, 1, 12, 24, 22, 15, 31, 18, 41, 75, 44, -5, -61, -73, 22, -41, -11, -3, 5, -5, 4, 50, 111, 86, 70, 67, 1, -9, -18, -30, -20, 7, 35, 33, 27, 13, 23, 27, 51, 54, 3, 8, 53, 27, -15, -27, -16, 44, -31, -33, 94, 89, 55, 14, -15, -12, 9, -13, -39, -24, -12, -18, 2, -10, -12, 2, 3, 11, 28, 24, 2, 32, -1, -13, -32, -33, -21, 4, 52, 66, 78, 43, 9, -6, 6, -1, -19, -36, -44, -31, -33, -31, -59, -32, -14, 14, 33, 53, -20, -10, -6, 16, -10, -21, -15, 11, 52, 84, 43, 33, 17, 34, 18, -22, -14, -54, -46, -17, -7, -24, -50, -65, -20, 28, 10, -10, -41, -57, -28, -18, -17, -17, 26, 99, 85, 85, 33, 26, 17, 25, -14, 11, -17, -64, -47, 29, 35, 15, -1, -24, -13, -9, 3, -26, -47, -13, -38, -16, 44, 8, 74, 77, 82, 63, 41, 16, 14, 9, -16, 22, 10, -8, 40, 86, 89, 84, 102, 58, -1, 4, -12, 0, -18, 1, -32, -9, 62, 65, 191, 94, 102, 36, -4, 2, -7, 9, 36, 45, 76, 49, 89, 103, 133, 119, 127, 60, 4, -22, -34, -32, -9, -28, -44, -17, 59, 82, 130, 78, 5, 14, -18, -34, -5, 16, 29, 44, 63, 75, 90, 75, 105, 135, 58, 53, -8, -74, -29, 39, 13, -29, -31, -25, 19, 38, 44, 8, 36, 22, -1, 0, -2, 25, 21, 24, 39, 33, 59, 52, 101, 80, 28, -17, -10, -41, -31, 16, -47, -66, -13, -36, 27, -6, -31, 46, 86, 55, 40, 31, 57, 5, 12, 12, 10, -3, 6, 34, 28, 35, 3, -18, -60, -26, 12, 0, -17, -59, 15, 9, -28, -64, -68, 121, 53, 55, 60, 52, 34, -45, -8, -44, -55, -79, -34, -25, 3, -21, -35, -43, -49, 45, 34, 20, -55, -28, -14, -22, -72, -72, -106, -3, -13, -5, 13, -24, -20, -51, -61, -67, -71, -107, -90, -71, -29, -25, -19, -6, 19, 90, 74, 17, -14, -58, 16, -43, -16, -47, -110, -9, -3, -23, -5, -28, -67, -55, -45, -104, -85, -72, -81, -3, 0, -39, -11, 11, 66, 60, 56, 51, 6, -19, -65, -28, -9, -9, -77, -16, -2, -48, 1, -18, -11, -32, -60, -45, -78, -54, -17, -4, -27, 9, -6, 11, 32, 0, 63, 8, 2, 14, -85, -7, -1, 15, -50, -7, 24, -33, -18, -6, -18, -28, -21, 11, -19, -24, -9, -34, 4, -1, 18, 37, 51, 49, 44, 13, 1, 28, -8, 11, 3, -3, -5, 50, -2, 39, 50, -7, -26, -2, 17, -1, 2, -13, 7, -18, 2, 24, 38, 79, 36, 21, 23, -8, -48, -26, -66, 7, 29, -43, 2, -19, 29, 45, 75, 25, 26, 16, 37, 24, 12, 24, 15, 12, 7, 23, 16, 27, 36, 17, -22, -69, -60, -57, -21, -13, 37, -8, 32, 13, -12, 7, 36, 53, 11, 41, 19, 24, 12, 29, 35, 71, 40, 49, 13, 13, -4, -45, -90, -33, -43, -34, -12, -19, 22, 4, 38, 1, 18, 36, -3, -29, -55, -33, 24, 9, -32, 11, -11, 18, 29, 38, 27, 4, 2, 13, -24, -47, -77, -18, -16, 5, 15, 14, 0, 9, 42, 25, 14, -49, -21, -3, -21, -16, -46, 18, 21, 2, 77, 36, 19, 14, -14, 17, -30, -48, -48, -18, -4, 20, -14, 20, -5, 44, 3, 30, 41, 7, -31, -52, -33, -58, -88, -12, -3, 56, 60, 71, 47, 50, 35, 34, 19, -4, 0, 16, 6, 1, -17, -20, 6, 6, -23, -23, -64, -53, -18, -10, 30, 54, -35, -23, 32, 9, 7, -15, -2, -8, -33, -24, 0, 6, -9, 1, -11, 20, -15, 2, -14, -5, 4, 18, 18, 9, 16, -16, -19, 19, 14, -15, -12, -22, -12, -20, -18, 7, -19, 11, -13, 19, 4, -11, -2, -11, 1103, 14, -3, 15, -19, -37, -36, -25, -44, -29, -33, -40, 3, 6, 30, -24, -3, -12, -31, -23, 11, 16, -4, -18, 5, 21, 19, -8, -10, 9, 6, -5, -3, 1, -42, -9, 36, -14, 28, 77, 52, 12, -9, 12, 45, 74, 15, -37, -11, -35, -26, -31, -6, -12, -3, -2, -11, -13, -2, 0, 50, 57, 7, 5, 67, 73, 83, 85, 60, 65, 20, 57, 33, 1, 47, -9, -35, -78, -71, -77, -84, -2, 11, 1, 9, 8, 8, 2, 72, 57, 11, 18, 89, 98, 87, 76, 76, 79, 24, 62, 52, 3, -5, 23, -21, -69, -79, -118, -107, -21, -17, 14, 6, -5, -9, 31, 16, 80, 114, 72, 109, 96, 68, 62, 102, 42, 59, 39, 0, -31, -30, -2, -16, -37, -70, -97, -7, 20, 11, -2, -10, -11, 2, 27, 28, 70, 100, 69, 60, 58, 82, 55, 37, 35, 29, 32, -3, -13, -55, 10, -34, -13, -29, -55, -18, 44, 9, 14, -11, -4, 24, 39, 14, 69, 106, 66, 66, 42, 32, 52, 13, 9, 23, 27, -16, -17, -40, 7, -9, -2, -7, -97, -62, -27, -18, -25, -12, -11, -45, 10, 41, 120, 153, 65, 10, 11, 21, -24, -12, 16, -5, -16, -7, -57, -27, -8, 2, 18, -29, -76, -98, -58, -6, -18, -18, -35, -60, 23, 87, 140, 80, -24, -6, -15, -48, -67, -41, -41, -2, 1, 17, -14, 26, 30, -9, -24, 4, -69, -79, -52, 2, -54, 15, -17, -93, -30, 45, 76, 13, -68, -59, -63, -95, -66, -57, -42, 3, 33, 32, 0, 42, 28, 20, -16, -2, -52, -45, 6, -58, 3, -1, 33, -48, 5, 22, 2, -63, -61, -69, -91, -75, -68, -38, -29, 2, 28, 18, 56, 49, 31, -4, -73, -43, -25, -22, -4, -54, -44, 20, -8, -3, 118, 3, -26, -54, -84, -130, -97, -83, -71, -41, -22, 33, 46, 43, 59, 53, -8, -41, -49, 1, -34, -20, -20, -37, -49, 6, 20, -51, 76, 38, -84, -126, -94, -101, -85, -52, -53, -31, 6, 35, 49, 43, 1, -19, -42, -47, -27, -11, -78, -61, -21, -73, -16, 29, 20, 2, 49, 9, -37, -89, -85, -58, -57, -25, -46, -13, 23, 37, 46, -11, 9, -51, -30, -37, -8, -26, -55, -38, -6, -95, -34, 10, 26, 8, 55, 31, -12, -56, -74, -34, 13, 6, -29, 4, -1, 23, 36, 13, -31, -27, -4, -1, 24, -26, -10, -26, 9, -102, -43, -5, -5, 54, 95, 71, -5, -54, -44, -41, 4, -14, -14, -44, -13, 58, 53, 13, -27, -11, 23, 8, 63, 46, 42, -2, 17, -64, -17, -34, 39, 123, 139, 92, 28, -73, -75, -61, -18, -9, -57, -61, -15, 87, 46, -23, -19, -10, 21, 37, 76, 56, 38, -20, -61, -108, -19, -18, 33, 111, 48, 63, 43, -44, -62, -29, -14, -15, -82, -88, -64, 38, 1, -15, 10, 42, 19, 69, 45, 40, -5, -19, -130, -81, -22, -14, 34, 76, 104, 32, -5, -28, -68, -33, -34, -53, -65, -66, -88, -7, -15, -2, 25, 46, 31, 23, 21, 5, -39, -109, -60, -72, -66, -9, 34, 13, 22, 58, 14, -5, -25, -58, -20, -62, -35, -40, -50, -21, 43, 26, 33, -2, -13, -8, -9, -32, -51, -121, -61, -59, -22, 33, -2, -12, 22, 18, -7, 3, 21, -30, -44, -42, -39, -21, 31, 25, 28, 1, 15, 25, -19, 5, -16, -42, -75, -97, -82, -22, -33, 16, -13, -21, 63, 26, -26, -2, -18, -4, 0, -51, -28, -21, 12, 40, 9, 55, 34, 27, -15, -13, -25, -85, -76, -124, -57, -28, -3, -10, 39, 73, 17, 1, -20, -1, 53, 75, 50, 16, 9, -17, 23, 16, 24, 10, 8, -4, -41, -46, -82, -77, -101, -81, -52, 18, 18, -15, 42, 69, 50, 45, 33, 2, 50, 53, 24, 4, 26, 16, 22, 21, -13, 5, 0, -17, -11, -51, -75, -96, -66, -50, -38, -46, 10, -6, 5, 12, 47, 53, 82, 63, 70, 5, 28, 80, 39, 3, 12, -6, 75, -1, -38, 23, 38, -18, -65, -38, -14, 12, 13, 9, -1, -2, -10, 19, 44, 35, 70, 48, 66, 82, 102, 80, 52, 51, 88, 69, 87, 94, 105, 98, 68, 59, 86, 43, 40, 9, -5, -1, -14, 9, 13, -2, -17, 17, 27, 53, 46, 79, 61, 94, 66, 18, 71, 16, 86, 93, 49, 55, 28, 10, 12, 29, 22, 11, -6, 13, 7, 17, -6, -10, 20, 4, -12, 1, 10, 9, 3, -9, -20, -4, 15, -1, 25, 11, 6, -3, 19, 8, 17, -11, 6, -14, 5, 11, 10, 17, -362, -10, -16, -3, -13, 5, -35, -28, -20, -15, 9, 33, 14, -31, 10, 29, 27, -1, 54, 39, 62, 51, 47, 26, -13, 15, 19, 5, 10, -11, 16, -12, -18, -52, -35, -86, -55, 22, 25, -8, 27, -4, -22, 11, 33, 4, -5, -52, -73, -22, -25, -43, -51, -11, 12, 12, -3, -12, 14, -1, 0, -32, -53, -105, -52, 51, -4, -1, -1, -28, -57, -27, -19, 11, -2, 12, 24, 4, 35, 36, 29, -17, 16, -13, -19, -18, -5, 14, 36, -95, -87, -106, -108, -70, -44, 4, 3, 3, 41, 20, 19, 6, -4, -21, -8, 31, 2, 29, 35, 57, 24, -16, -13, -8, -38, 2, 14, -65, -88, -97, -112, -65, -36, 10, 4, 14, -5, 48, 26, 40, 25, 38, 45, 60, 51, 25, -4, 8, 42, 13, 18, 10, -21, -36, -42, -26, -38, -84, -124, -55, -35, -23, -27, -5, -6, 23, 27, 32, 9, 25, 43, 76, 33, 21, -49, 11, 59, 23, 15, -1, 26, 27, -35, -39, -46, -73, -53, -1, -18, -10, -29, 5, -21, -10, 26, 23, 49, 27, 50, 53, 41, -20, 14, 17, 39, 18, -6, 10, 19, -35, -14, -10, -13, -40, -6, 1, 2, -26, -11, -46, -23, 1, 34, 63, 90, 75, 74, 58, 58, 31, 19, 6, -11, 12, 10, 4, 54, 14, 15, 33, 12, 17, 16, -25, 6, 28, -33, -56, -55, 13, 53, 66, 90, 57, 31, 26, 20, 1, 4, -16, -1, 65, 21, 19, 11, 40, 23, 51, 16, -2, -37, -44, -28, 7, -16, -48, -75, -12, 40, 80, 75, 15, -5, -14, 1, -23, -14, -1, -1, -7, 49, 48, 91, 27, 31, 38, 22, 11, -22, -7, -63, -5, -33, -46, -78, 3, 75, 88, 33, 14, -38, -9, -33, 6, -7, 2, -25, 28, -17, 38, 93, 24, 35, 49, 28, 0, 23, 8, -21, -41, -31, -58, -16, 46, 107, 55, 36, -22, -34, -44, -22, 8, -3, -8, 14, 37, 4, 36, 44, 35, 71, 38, -5, 32, 21, -3, -17, -49, -66, -39, 23, 78, 61, 34, -6, -17, -51, -40, -46, -12, -38, -69, 5, 8, -10, 45, 92, 61, 65, 14, 14, 11, 14, 14, 1, -39, -76, -38, 16, 32, 14, -24, -58, -44, -58, -40, -52, -38, -87, -101, 15, -7, 12, 53, 87, 59, 39, 27, 26, 7, -14, -4, -9, -46, -73, -69, -11, 14, -9, -69, -86, -61, -68, -68, -75, -75, -129, -29, 48, 24, 7, 11, 56, 88, 52, 21, 38, 20, 3, 3, -24, -40, -57, -25, 58, 4, -45, -75, -51, -23, -34, -30, -31, -79, -74, 4, 5, 25, -21, 19, 68, 79, 104, 50, 16, 62, 39, -10, 17, 18, 26, 53, 93, 29, -16, -7, -39, -33, -21, 3, -10, -43, -9, 66, 49, 65, 16, 39, 47, 15, 63, 76, 56, 55, 46, 29, 77, 96, 107, 74, 108, 66, 41, 39, 29, 26, 12, -1, 12, 7, -2, 109, 84, -11, 21, -8, 24, 32, 16, 59, 55, 72, 32, 54, 41, 89, 84, 64, 54, 40, 14, 5, 38, 1, 8, 36, 2, 46, 26, 96, 85, 43, 18, 52, -11, -87, -3, 76, 59, 37, 2, 11, 25, 43, 40, -1, 13, -4, 27, -15, 14, -1, 19, 39, -12, -2, 26, 76, 24, 20, 49, 5, -42, -6, -45, 25, 11, 14, -17, -42, 8, -2, -37, -27, -24, -33, -22, 4, 22, 35, 38, 18, 15, 46, 34, 35, 16, 37, 14, 23, 2, -60, -71, -43, 2, 33, -30, -43, -3, -28, -7, -9, -35, 9, -8, -12, 25, 32, 32, 18, 39, 5, 11, 67, 16, 13, -12, 7, 48, 13, -40, -35, -4, 18, -16, -29, -25, -24, -11, 14, -1, -1, -17, 16, 0, 37, 39, 32, 3, -5, 20, 28, -15, 19, 10, 13, 58, -22, -64, -53, -38, -57, -32, -26, 10, -3, 28, 32, 29, 14, 24, 69, 34, 36, 54, 14, -41, -27, -13, 61, 11, 11, -5, -1, 16, 24, -19, -35, -56, -52, -6, -21, 9, 6, 17, -13, 5, 12, 55, 62, 39, 17, 15, -13, -42, 3, 3, 34, 16, -11, -19, 9, 10, 21, 0, 1, -26, -17, -19, -49, -3, -27, 6, -56, -104, -53, -13, -28, -9, -5, -56, 2, -36, -17, 34, 38, 9, -3, 0, -2, -16, 4, 0, 35, 10, -32, -13, -12, -51, 22, 50, 46, -25, 11, 9, 33, -68, -16, -36, -20, 11, -13, 13, -10, -2, 14, 11, -17, -7, -3, -11, 7, 2, -10, -6, 17, -21, -8, 2, 5, 12, -26, -11, -9, -19, -2, 12, 2, 13, -13, 6, -7, 2, -19, -1, 692, 15, 17, -13, -8, 0, -32, -17, -44, -10, 2, -13, 10, 20, -17, -29, 0, -11, -43, -33, -40, -43, -9, 5, -5, -2, 15, -13, -11, -4, -10, -22, 0, 37, -4, -4, 19, -28, -12, 30, -4, -13, -65, -53, -13, -18, -43, -18, -63, -59, -65, -33, 69, -6, -7, -11, 19, -6, -15, -23, -6, 15, 39, 41, 47, 26, 19, 59, 4, -19, -23, -32, -12, -1, -30, -61, -64, -79, -68, -134, -77, -14, -1, 11, 15, 15, -9, -8, -19, -2, 6, -6, 25, 20, 20, -12, 37, 26, 25, -1, -8, -3, -16, 0, 2, -25, -55, -71, -82, -58, -33, 7, 18, 16, -17, -37, -89, -42, -46, -15, -33, -9, -14, 2, 25, 12, 54, 5, 28, 15, -3, -13, -6, -25, 0, -24, -33, -13, -37, -2, 3, -14, -13, -22, -20, -25, -67, -97, -40, -17, 6, 31, -18, -16, 11, -11, 13, 18, -5, 9, -33, -34, -45, -54, -41, -20, -66, 15, 0, 2, -7, -48, -33, -61, -86, -56, 0, -11, -25, 21, -50, -24, -60, -34, -3, 16, -6, -1, -16, -43, -30, -70, -87, -108, -34, -27, 1, 30, -6, -59, -70, -43, -108, -97, -23, 1, -20, 18, -7, -36, -40, -61, -4, 48, 14, -35, -43, -74, -44, -64, -97, -123, -37, -3, -19, 5, -24, -81, -78, -79, -118, -112, -11, -10, -9, -14, -21, -21, -3, -20, 0, 1, -24, -9, -18, -43, -47, -60, -46, -57, -59, -42, -16, 15, -14, -72, -97, -126, -109, -97, -18, -27, -34, 8, -33, 7, 32, 14, 0, 6, -4, 10, 13, 18, 21, -3, -11, -67, -43, -7, -43, -69, -42, -119, -108, -101, -98, -71, -45, -38, -9, -3, -39, 21, 14, 3, -16, -9, -6, -10, -59, -35, -8, 4, 17, -12, -48, -50, -11, -35, -98, -111, -138, -135, -109, -101, -54, -33, -15, -26, -26, 3, 41, 20, -21, -46, -62, -66, -90, -81, -29, -9, -48, -3, -39, -27, 2, -38, -102, -123, -145, -155, -104, -59, -37, -23, -40, -35, -34, -16, 59, 12, -17, -44, -18, -69, -56, -82, -39, -39, -33, -8, -1, -25, 35, -35, -80, -111, -150, -173, -149, -95, -19, -28, -65, -30, 8, 7, 76, 40, 19, 31, -7, -21, -44, -82, -79, -28, -71, -32, -31, -12, 16, -40, -65, -103, -112, -160, -144, -97, -14, -45, -73, -43, 11, 33, 65, 62, 81, 82, 11, 18, -54, -80, -87, -52, -95, -48, -73, -26, -1, -35, 41, -29, -28, -56, -55, -65, -48, -91, -103, -37, 0, 6, 23, 54, 79, 73, 52, 2, -62, -83, -79, -93, -59, -31, -18, -23, 6, -30, 58, 76, 119, 86, 2, -39, -102, -88, -111, -104, -67, -50, -10, 19, 87, 69, 26, -13, -61, -88, -98, -72, -86, -82, -6, -22, -6, -37, 67, 96, 102, 63, 9, -9, -34, -53, -68, -64, -88, -64, -30, -5, 72, 57, 42, 10, -32, -72, -98, -98, -46, -91, -62, -20, -9, -26, 33, 74, 126, 56, 35, 49, 5, -12, -11, -8, -10, -54, -53, 7, 17, 77, 3, -16, -52, -75, -72, -83, -52, -104, -67, -61, -5, -4, 17, 89, 85, 76, 23, 50, 30, 40, 31, 9, -34, -36, -32, 2, 55, 60, -5, -17, -50, -38, -45, -43, -77, -70, -63, -71, -25, -15, -1, 14, 31, 46, 80, 50, 52, 61, 34, -32, -37, -3, -16, 4, 2, 49, 24, -21, -62, -86, -132, -73, -73, -88, -42, -37, -7, -7, 42, 89, 36, 52, 41, 5, 76, 43, 9, -21, -54, -52, -14, -19, -7, -18, -27, -51, -90, -116, -161, -101, -89, -46, -20, -26, -3, 17, 37, 33, 0, 0, 19, -28, 31, -12, -18, -6, -40, -45, -21, -36, -38, -32, -52, -50, -100, -149, -115, -73, -46, -36, -8, 19, 12, -19, 37, 47, 37, 55, -8, -45, -29, -72, -59, -20, -32, -45, -19, -38, -42, -40, -33, -38, -122, -94, -77, -74, -36, -52, -24, 3, -12, 2, 4, -36, -45, -22, 18, 1, -73, -88, -92, -95, -90, -55, -53, -86, -40, -111, -91, -67, -78, -22, -25, -19, -24, -33, 0, 10, -12, 2, 3, -20, -33, -69, -31, -27, -13, 25, -32, -22, -28, -48, -3, 39, -2, -51, -79, -58, -43, 1, -25, 1, -21, -2, 13, -3, 3, -1, 13, 12, -21, 11, -6, 18, 13, 7, 15, -30, -40, 3, 37, 8, 17, -8, 21, 8, 12, 4, 5, -18, 20, -16, 20, 19, 2, 18, 3, -16, -3, -15, 9, -4, -3, -12, -7, 9, 4, -19, 5, 14, -2, -18, 4, -10, 15, -14, -6, -19, 9, 4, -10, -3, -1, 228, 13, 7, -20, -12, -7, -60, -75, -38, -66, -40, -38, -73, -54, -65, -54, -69, -27, 31, -56, -3, -29, -19, -14, 8, 1, -13, -11, 2, 9, -4, -18, 9, -45, -50, -74, -44, -7, -40, -11, -47, -76, -97, -61, -53, -52, -50, -124, -97, -41, -23, -29, -20, 11, 11, 17, 12, 1, 6, 24, -28, -93, -100, -62, -2, 2, -8, 31, -8, -16, -48, -47, -64, -29, -57, -42, 1, 29, 50, 36, 36, 4, -9, -16, -10, -17, 10, 25, 40, -50, -25, 14, -28, -13, 10, 5, 23, 27, 10, -12, 26, -35, -47, 9, 70, 45, 48, 16, 23, 2, -27, -15, -7, -16, -24, -18, -2, 0, 7, -6, -24, -29, -33, -28, -22, -14, -49, -13, 27, 61, 62, 67, 106, 93, 26, -6, -37, -7, 21, 8, 4, 14, -6, -7, -17, -8, 45, -24, -67, -47, -46, -42, -87, -85, -77, -42, -4, 42, 47, 106, 95, 77, 57, 1, -43, 19, 54, -18, -5, -8, 31, -18, -21, 21, 25, -13, -58, -48, -71, -83, -77, -75, -69, -24, 19, 43, 65, 58, 18, 28, -3, -56, -44, 25, 40, 33, -15, -5, 41, 12, -9, 12, -12, -6, -35, -67, -51, -40, -58, -50, -78, 31, 96, 113, 77, 23, 15, 40, -6, -22, -10, 0, -26, -5, -17, 4, 66, 35, 24, 23, 14, -39, -65, -53, -36, 12, -41, -37, -81, 39, 105, 73, 70, 12, -17, -12, -27, 2, -3, -35, 4, 27, 8, 40, 67, 65, 56, 48, 3, -55, -56, -41, -18, -9, -1, -32, -47, 27, 95, 58, 28, 10, -1, 6, -18, 7, -9, 0, -8, -15, 45, 58, 76, 74, 47, 7, -7, -14, -62, -42, -30, -5, 38, -14, -23, 93, 136, 71, 38, -27, -38, -10, -21, 12, 24, 26, -3, -26, 14, 66, 86, 34, 62, 28, -17, -22, -53, -43, -20, 33, 34, 9, 42, 112, 102, 74, 12, -47, -61, -16, 3, -7, 46, 33, -18, -24, 17, 39, 48, 35, 61, 20, 0, -36, -55, -21, 21, -15, -5, 21, 82, 110, 92, 50, -49, -52, -74, -48, -10, 16, 18, -38, -45, -37, -3, 23, 97, 46, 37, 3, -32, -15, -58, -34, -18, -43, -44, 6, 86, 120, 97, 43, -19, -60, -38, -11, -1, -19, -43, -48, -50, -33, -1, 42, 74, 59, 39, -13, -12, -19, -45, 1, -26, -60, -65, -54, 30, 115, 65, 27, -30, -30, -26, -47, -23, -69, -85, -70, -2, -4, 17, 15, 36, 77, 76, -1, 0, 5, -16, 6, -31, -68, -86, -73, 49, 51, 12, -53, -37, -32, -42, -8, -33, -41, -66, -70, -36, -21, -12, 7, 87, 92, 94, 68, 20, 18, 5, -15, -21, -53, -91, -30, 58, 30, -44, -27, -42, -23, 11, -6, 23, -31, -54, -42, -34, 16, 2, 35, 66, 15, 51, 74, 60, 47, 54, 6, 28, 1, 32, 23, 56, -9, -43, -21, 7, -16, 4, 2, -3, 14, -21, -3, -29, -39, 2, -8, 45, 47, 66, 81, 81, 41, 39, 49, 39, 54, 62, 37, 30, 0, -31, -13, 11, -18, -31, -17, -44, -8, -20, 3, -21, 19, 17, 41, 25, 18, 57, 81, 66, 1, 39, 46, 29, 64, 75, 22, 12, -15, -6, -24, 29, 15, -48, -35, -21, -33, -21, -65, -25, 24, 24, 45, -42, 6, 37, 75, 57, 29, 21, 13, 30, 23, 6, 2, -24, -23, -5, -2, -6, -11, -36, -45, -10, -28, -16, -66, -23, 52, 5, 14, -19, 1, 45, 63, 75, 29, -23, 15, 20, 44, 23, -5, -27, 6, -15, -36, -11, -30, -53, -34, -53, -54, -38, -50, -45, -5, 5, -26, 45, 3, -32, -13, 2, 8, -18, 13, 25, 30, 39, -22, -17, -28, -54, -27, -47, -48, -45, -43, -31, -55, -23, -13, -12, -10, 16, 39, 65, 15, -82, -72, -75, -95, -48, -17, -3, 58, 18, -6, -31, -31, -42, 19, -27, -29, -27, -15, -24, -10, -51, -20, 20, 12, -17, -20, -19, -35, -36, -54, -33, -54, 24, 10, 32, 8, 27, -11, -32, -35, -3, 18, 21, 33, -17, -32, -28, -2, -24, 14, 10, 8, 20, -6, 10, 3, -3, 11, -35, 1, -13, -12, -20, -21, -11, -17, -61, -12, -16, 8, 24, 6, 8, -11, -7, -9, 10, 45, -5, -2, 11, -15, -15, -16, -7, 38, -6, -29, -45, -8, -29, 26, 42, 33, -38, 26, 2, 32, -22, -24, -6, -25, 2, 16, -4, -15, 9, -13, -15, 16, 11, 7, 13, -3, 0, 2, -13, 0, 1, 17, -18, 10, 12, -20, -12, -6, 6, -12, 15, -14, -9, -10, -8, -19, -19, -19, 2, 1180, -2, 4, -18, -4, -48, 0, -5, 17, -7, -2, -48, -54, -33, -32, -124, 8, 2, -10, -12, 4, 2, 9, -29, -18, -15, 20, 3, 12, -10, 4, -4, -2, -13, -11, 26, 70, 110, 65, 6, 39, 27, 33, 36, 77, 78, 58, 40, 35, 39, 64, 35, 37, 26, -6, -18, 9, -21, -4, -8, 50, 41, 76, 91, 89, 126, 88, 61, 19, -13, 4, 53, -8, 7, 41, -2, -6, 23, 22, -4, -30, -20, 27, 8, -14, -9, -21, -55, 41, 64, 31, -1, 40, 75, 87, 48, 12, 24, 18, 46, 28, 43, 26, 5, 6, -4, -16, 7, 45, 73, -13, 6, -6, -19, 26, 1, 9, 25, -5, -34, -6, -20, 5, 28, 11, 21, 40, 33, 4, -2, -20, -7, -20, -48, 6, -1, 76, 95, 27, -5, 3, 7, 29, 44, -31, -27, -81, -52, 0, -38, -2, 20, 30, 27, 38, 23, 6, -41, -31, -39, -38, -37, -6, -51, 2, 40, -8, 2, 11, -21, 37, 25, -56, -56, -38, -55, 1, -21, -6, 14, 24, 40, 64, 34, 15, -1, -45, -42, -30, -1, -1, -37, -25, -8, -11, -2, -12, -6, -52, 35, -1, 1, -20, -3, -6, -11, 0, -9, 3, 20, 34, 46, -6, -15, -46, -31, -52, -28, -25, -14, -44, 21, 31, -7, 15, 10, -27, -22, 53, 30, 4, -7, 6, 10, -3, -3, -1, 24, 42, 51, 41, 12, -12, -43, -18, -65, -45, -20, -39, -40, 48, -9, 8, -13, -8, 25, 71, 46, -11, -31, -24, -7, -12, 22, 23, 27, 38, 39, 17, -1, 48, -10, -6, -17, 28, -11, -33, -4, 2, -16, 33, 4, -65, 12, 36, 30, -16, -55, -5, -25, -34, -2, 20, 28, 37, 26, 17, 28, 52, 33, 11, 5, 28, 16, -48, 26, -31, 16, 14, -6, -3, 52, 54, 59, -7, -28, -39, -51, -12, -11, 37, 3, 30, 10, 25, 62, 58, 25, -13, 7, 21, -4, 3, -7, 10, 2, -31, -29, -49, 68, 81, 29, -18, -23, -14, -26, -13, 6, -3, 47, 37, 18, 53, 60, 20, 16, -21, 12, -40, -36, -48, -28, -43, 29, 0, -35, -27, -17, 30, 80, 29, -3, -18, -23, 24, -20, 15, 55, 50, 47, 59, 35, 3, -26, -36, -10, -47, -64, -60, -27, -90, -36, 29, -35, -30, 12, 39, 104, 23, 3, 35, 42, -4, -27, -8, 45, 82, 125, 60, 17, 14, -4, -40, -5, -42, -28, -5, -9, -66, -40, -8, -12, 18, 36, 32, 91, 0, -25, -10, 16, -31, -72, -5, 74, 136, 120, 48, 1, -40, -5, -20, -3, -21, -25, -10, -22, -48, -71, -5, 23, 76, 85, 81, 44, -18, -31, 1, -48, -97, -80, -25, 100, 179, 128, 20, -18, -53, -22, -17, -3, 0, -15, 46, -55, -37, -64, -17, -12, 89, 90, 90, -4, -49, -66, -72, -82, -120, -129, 14, 183, 229, 128, 17, -5, -34, -11, -29, -34, 8, -43, 27, -24, -59, -72, -34, 15, 99, 82, 44, -28, -53, -58, -97, -100, -120, -98, 28, 198, 170, 84, 2, -31, -27, -41, -19, -15, -22, -38, -15, -22, -10, -66, -22, 38, 29, 20, 34, -44, -78, -48, -68, -98, -166, -65, 84, 143, 109, 23, -29, -22, -32, -37, -28, -33, -3, 30, 14, -52, -72, -22, 12, 18, 8, 36, 15, -59, -85, -63, -124, -126, -113, -53, 91, 146, 80, -12, -39, -39, 19, 34, 32, 24, -6, 38, -25, -105, -27, -10, 0, 30, 24, 45, 40, -52, -60, -60, -92, -90, -77, -16, 62, 101, 102, 30, -10, 39, 18, 8, 36, 40, 5, -1, 20, -73, 2, 3, -19, 52, 87, 55, -2, -35, -18, -23, -57, -79, -40, -18, -1, 62, 58, 66, 42, 41, 37, 29, 23, 7, 13, -19, 15, -52, 21, -1, 12, 72, 79, 76, 34, 15, -27, 9, -56, -41, -32, -50, -7, 27, -10, 15, 50, 41, 43, 36, 44, 33, 52, 35, 47, -15, -2, 0, 0, -4, 41, -2, 34, 88, 60, 33, -6, 11, -30, -89, -63, -31, -33, 41, 133, 57, 84, 104, 84, 61, 62, 39, 29, 37, -6, 1, 17, -18, -14, -6, 34, 53, 48, 39, 5, -2, 4, -28, -25, -7, 1, 25, 140, 143, 116, 96, 76, 67, 42, 29, 36, 21, 6, -4, 12, -13, -20, 17, 11, 45, 32, 37, 31, 31, 56, 64, 5, 12, 8, 24, 62, 56, 69, 36, 36, 48, 44, 30, -10, -20, 2, 5, -18, 0, -7, 7, -20, 9, 16, 18, -3, -6, 5, 17, 21, 3, -24, 10, 12, 2, -10, 6, 13, -2, 18, -8, 15, 13, -9, -15, 20, 126, -13, -5, -9, -19, -1, -22, -16, -49, -63, -69, -87, -72, -102, -131, -110, -80, -46, -37, -37, -26, -21, -17, -22, -23, 17, -8, -12, -16, -17, 20, -2, -4, -53, -83, -85, -99, -119, -153, -117, -117, -121, -213, -148, -158, -80, -101, -124, -112, -117, -78, -64, -58, -22, 12, 4, -19, -2, 44, 20, -24, -34, -36, -34, -26, -74, -80, -44, -47, -15, -57, -97, -109, -55, -120, -122, -100, -68, -43, -100, -86, 9, -7, 9, -6, -2, 15, 24, -12, -58, -33, 47, 8, -17, -5, -42, -44, -48, -75, -68, -63, -78, -109, -85, -81, -27, -37, -50, -56, -29, -2, -14, -14, -13, 30, -28, -77, -63, -35, 7, -11, -24, -45, -82, -65, -44, -58, -63, -77, -92, -102, -86, -73, -36, -4, -6, -20, -23, 11, -8, -3, 0, 49, -20, -50, -61, -13, -13, -29, -56, -52, -78, -42, -47, -75, -83, -84, -88, -44, -58, -91, -45, -54, -6, 3, 26, -30, 6, 8, 11, 75, -19, -25, -49, -36, -17, -73, -63, -24, -33, -45, -50, -39, -11, -40, -63, -43, -52, -34, -64, -66, 7, 36, 35, -34, -6, 19, -13, 38, -39, -31, -65, -55, -17, -30, -45, 24, -7, -11, -5, -4, 13, 28, 31, 0, -21, -29, -33, -84, -31, 13, 35, -15, -53, -3, 44, 7, 31, -5, -16, -29, -14, -23, -59, 46, 53, 52, 28, 42, 14, 41, 48, 25, 5, 7, -29, -55, 0, 9, 49, -20, -24, -5, 31, -21, 38, 32, -11, -27, -21, -24, -21, 21, 50, 70, 36, 60, 36, 54, 10, -23, 34, 8, 10, 9, -1, 23, -9, -35, -22, -16, 19, -27, 51, -52, -35, 6, 33, -10, 5, 43, 49, 47, 63, 49, 0, 2, -8, 18, 5, 8, 0, 43, 37, 15, -6, 6, -12, 4, 24, 40, 93, 16, 15, 8, 20, 28, 15, 30, 45, 61, 45, 67, 44, 3, 15, -1, -17, -10, 28, 45, 0, 3, 37, -1, -33, -1, 34, -3, 40, 17, 14, 21, -11, -9, 37, 9, 43, 47, 46, 46, 53, 55, 51, 17, -1, 29, 51, 27, 44, 43, 76, 36, -2, -7, 0, 8, -4, 48, 55, 49, -7, 6, 29, 13, 38, 45, 18, 55, 39, 52, 34, 43, 39, 42, 42, 53, 63, 9, 31, 16, 0, 27, 26, -1, 2, 29, 56, 47, 48, 5, 40, -2, 20, 13, 44, 7, 58, 70, 4, 42, 37, 50, -10, 21, 45, -33, -32, -38, -26, -12, -15, -13, -10, -25, -13, 1, 10, 26, 16, -38, -32, 26, 22, 28, 17, -13, -18, -19, -8, 35, 11, -34, -19, -51, -14, -32, -1, 8, -20, -83, -74, -53, -55, -4, 30, 3, -21, -58, -49, 13, 13, 10, -62, -71, -80, -45, -1, 0, -3, -4, 16, -32, -4, 0, 6, -14, -30, -73, -16, 2, -12, 10, 41, -7, -60, -36, 8, 2, 12, -29, -70, -109, -90, -51, -37, -7, -4, -20, 4, -5, -44, -18, -8, 3, 14, -36, -63, 2, -39, -32, -7, 3, -61, -43, -24, 12, 11, -32, -50, -78, -90, -49, -48, -38, -24, -51, -2, -33, -13, -4, -27, 12, -51, -22, 30, -32, -25, -48, -25, -32, -97, -61, -20, -54, -1, -26, -67, -104, -99, -39, -23, -39, -20, 17, -3, 7, -16, 10, -19, 24, -11, 32, 51, 25, -38, -19, -59, -63, -88, -76, -41, -34, -15, -39, -139, -125, -95, -69, -44, -23, -36, 0, 22, 45, -30, -27, -20, -3, 5, 33, 1, 0, 27, -3, -55, -74, -102, -64, -31, -33, -21, -42, -133, -151, -118, -96, -34, -1, -23, 12, 35, 22, -40, -13, 12, 16, 47, 28, -7, 39, 21, -42, -54, -55, -54, -64, -34, -39, -2, -14, -68, -92, -69, 7, 1, 60, -6, 27, 17, 56, -25, 1, -7, 17, 17, -36, -53, 5, 29, -10, -3, -9, -39, -59, -58, -65, -49, -12, -9, 13, 15, 53, 63, 73, 30, 46, 21, 5, -69, -16, -14, 13, 20, 21, -27, 20, 17, -2, 31, 18, -16, -67, -49, -33, -10, 4, 1, 6, 63, 66, 109, 53, 16, 49, 24, 23, -33, -16, 14, 19, -1, 13, -18, 10, 35, 41, 52, 26, 2, -7, 26, 4, 9, 41, 41, 95, 120, 78, 65, 59, 10, 13, 28, -28, -10, -7, -19, 16, -13, 9, -5, 2, 30, 43, 40, 28, 46, 60, 34, 21, -41, -64, -14, 13, 19, 14, 12, 36, 26, 29, -9, 4, 14, 8, 21, 8, -8, -15, -1, -12, 11, -1, -2, 10, 12, 9, -12, -14, -20, -19, 12, 12, -15, -9, -3, 9, -19, -8, 17, 19, 6, 8, -4, 15, -961, 1, -15, -10, 0, -53, -25, -31, 5, -6, -33, -38, -48, -41, -33, -75, -20, -26, -45, -65, -63, -46, -56, -16, -8, 1, -6, 7, -4, -13, -11, -15, -8, -4, -36, -35, -70, -91, -98, -121, -67, -67, -73, -56, -15, -49, -111, -83, -20, 11, 70, 57, 68, 7, 5, 19, 20, 17, 31, 47, -38, -58, -73, -80, -121, -130, -128, -137, -63, -41, -57, -85, -103, -68, -74, -98, -21, 25, 26, -26, -35, -23, 17, 14, -17, -5, 39, 54, -5, -63, -109, -80, -130, -125, -61, -49, 8, 24, -4, 36, 46, 70, 36, 30, -3, -5, -44, -52, -51, -56, -25, 5, -11, 7, -65, -46, -40, -59, -45, -65, -76, -18, -32, -43, 17, 7, 22, 38, 28, 30, 15, 44, 46, 25, 3, -27, -108, -32, -21, -9, -9, -5, -27, -59, -38, -80, -28, 4, -30, -20, -26, -58, -30, -1, -2, 24, 29, 3, 31, 14, 13, 6, 38, 3, -36, 37, 32, -15, -5, 22, 29, -51, -21, -33, 5, 11, -11, -23, -15, -42, -54, -15, -27, -32, -12, -10, -19, 10, 5, 0, 30, -5, 5, 31, 49, 8, -1, -15, 1, -37, -24, 4, 8, 38, -3, 21, -36, -46, -55, -21, -43, -77, -18, -10, 35, 25, -4, 36, -2, 9, 11, 12, 26, 6, 14, 10, -1, -46, -13, 14, 68, 39, 15, -1, -34, -52, -18, -38, -65, -67, -56, -8, 44, 65, 41, 46, 21, -20, -2, 2, -42, -34, 5, 25, -18, 65, 9, 20, 40, 31, 11, -27, -9, -63, -32, -4, -51, -60, -32, -16, 84, 71, 50, 42, 21, 17, -4, -45, -37, -6, -24, 68, -2, 118, -6, -12, 45, 21, 22, 5, -24, -33, 22, 18, 1, -28, -5, 67, 116, 68, 60, 54, 44, 11, -32, -44, 16, -36, -3, 25, 21, 54, -41, -21, 24, 39, 10, -12, -9, -12, 3, -3, -3, -69, 13, 92, 80, 85, 99, 97, 97, 42, -1, -4, 14, -26, 9, 16, -16, 7, -11, 31, 51, 48, 37, 11, -23, -15, -19, -55, -43, -43, 33, 51, 72, 57, 92, 126, 81, 80, 42, -3, 4, -3, -15, 45, 33, 50, 55, 61, 63, 52, 3, 2, 5, -21, -22, -53, -38, -20, 31, 72, 38, 56, 48, 65, 65, 94, 25, -4, -10, 24, -33, 41, 10, 44, 126, 123, 109, 47, 11, 9, -1, -19, 0, -11, -12, -1, 32, 26, -9, -21, 8, 27, 55, 18, -18, -7, -31, 8, -11, 0, -77, -2, 173, 144, 124, 46, 15, -5, -13, -16, -49, -56, -32, 27, 22, -20, -57, 12, -21, -19, 24, 33, -19, -3, 26, 14, 8, -44, -74, -65, 66, 84, 41, 62, 29, 15, -67, -38, -76, -94, -20, 0, -20, -63, -35, 18, -47, -23, 4, -10, -37, 4, 10, 16, 1, -60, -112, -172, -22, 14, 45, 44, 35, 11, -1, -16, -73, -50, -7, 36, -6, -18, -21, -25, -47, -35, -45, -5, -28, 13, -20, -15, -33, -55, -142, -152, -49, 6, -47, 20, 60, 39, -42, -49, -43, -44, -20, 26, -9, -42, -13, -10, -51, -80, -90, -111, -13, -6, -2, -66, -4, -59, -54, -123, -60, -20, 4, 0, 20, -6, -15, -11, -7, -45, -15, 21, 6, 4, -35, -44, -68, -103, -71, -64, -4, 4, -3, -7, 51, 15, -35, -45, 20, -13, 37, 16, -22, 11, 17, 17, -37, -8, -15, 8, -1, -37, -26, -84, -119, -103, -74, -71, -29, -49, 15, -50, -18, 2, -56, -21, -28, 10, 42, 24, -30, -27, 7, -16, -8, -36, -20, -12, -36, -48, -75, -109, -103, -85, -70, -25, -4, -31, -18, -27, -12, 19, -16, -9, -10, -42, -25, -9, -45, -8, -1, 9, 27, -2, 19, -14, -33, -50, -47, -69, -19, -27, -13, -63, -10, -36, -18, 9, -3, 17, -8, -37, -31, -4, 5, -13, -43, -37, -67, 5, -3, 6, -22, -1, -6, -19, -20, -12, 9, 4, 13, -13, -10, -43, -35, 15, -15, 11, 29, -6, 10, 37, 7, 4, -36, -24, -8, -3, 34, 13, 81, 56, 6, 72, 37, 29, 12, 12, -14, 0, 2, -9, -23, 10, 18, 16, -19, -23, 22, 11, 41, 59, 27, 3, -43, -42, 5, 24, 71, 81, 75, 71, 73, 50, 108, 118, 74, 29, 15, 16, -18, 17, -11, -1, -15, -4, 16, 29, 55, 67, 86, 60, 74, 57, 38, 7, -21, 138, 84, 81, 55, 51, 41, 55, 55, 5, -10, 13, -18, 4, 7, -7, 11, -5, -14, 0, 18, 12, 8, -9, -17, 9, -10, 0, 1, 4, 14, 10, 11, 17, -13, -9, -4, -20, 6, -16, -12, 16, 16, 277, 2, 14, -2, 6, 37, -13, 12, -3, -31, 7, 28, 28, -9, 6, 58, 0, 0, 25, 11, -32, -17, 10, 20, 29, 6, -17, -2, -10, -13, 15, 15, -21, -15, 19, -8, -59, -35, -39, -9, 5, 34, -19, -24, -41, 55, 50, 28, 9, -1, -68, -37, -70, -17, -7, -11, -16, -11, -35, -13, -17, 19, -15, -5, -50, -39, -40, -22, -4, 53, 26, 54, 107, 110, 111, 143, 168, 101, 36, 12, 70, 47, 2, 10, -20, -4, -21, -36, -49, -34, -75, -100, -47, -24, -28, -42, 7, 36, 50, 53, 75, 92, 74, 30, 43, 98, 92, 88, 73, 79, 68, -6, 7, -4, 3, -46, -86, -142, -115, -76, -33, -28, -47, -13, 1, 18, 25, 3, 22, 15, 30, 1, 12, 30, 36, -7, 42, 12, 13, 0, 18, 7, -18, -55, -122, -112, -88, -100, -51, -16, -77, -27, -12, 8, -20, -5, -17, 19, -3, 4, -3, 1, -4, -14, 2, -20, -42, -4, 19, -13, -45, -74, -123, -114, -91, -78, -52, -59, -59, -45, -42, 25, -24, 4, 4, -37, -51, -11, 3, 7, 16, -38, -23, -39, -29, 4, 10, 20, -3, -96, -100, -114, -118, -79, -71, -77, -46, -3, 12, 2, 12, -20, -40, -41, -41, -3, 10, -12, -18, -25, -44, -2, 2, 22, 2, -14, -26, -52, -69, -140, -149, -51, -31, -46, -17, 8, 16, 58, 52, -6, -39, -49, -19, 2, -15, -4, -12, 26, -20, 4, 25, 35, -11, -57, 34, -73, -82, -74, -63, -27, 29, -9, -4, 22, 43, 58, 55, 27, -11, -27, -60, 0, -36, -28, -1, 0, -5, 14, 67, -6, -17, -43, -23, -104, -20, -2, -19, -20, -21, -31, 17, 60, 85, 61, 58, 21, -21, -46, -27, -19, -5, -11, -18, -21, 6, -14, 40, 20, -15, -82, -87, -120, -49, -54, -19, -10, 15, -2, 5, 7, 60, 40, -12, 18, -14, -15, -10, 23, 2, -22, -37, -63, -36, 18, 48, 28, -18, -46, -47, -94, -73, -26, -37, -62, -34, -18, -7, 50, 28, -8, -8, 24, 29, 19, 23, -8, -6, -18, -21, -63, 2, 23, 75, 45, 9, -35, -102, -56, -74, -54, -69, -50, -33, -15, -6, 24, 9, -20, -18, 5, 9, 3, 9, -5, -9, -42, -58, -34, 18, 55, 68, 43, 12, -64, -34, -22, -101, -135, -83, -23, -27, -26, 0, 4, -1, 4, 23, 38, 25, 61, 10, 16, -21, -35, -56, -61, -13, 35, 75, 48, 6, 4, 11, -25, -69, -101, -65, -36, -36, -13, 13, -13, 53, 58, 100, 72, 57, 64, 41, -4, -39, -15, -66, -27, -21, 27, 45, 51, 36, 35, 83, 74, 16, -19, -30, -46, -13, -3, 7, 26, 35, 105, 102, 66, 62, 21, -1, -22, -56, -28, -53, -39, 43, 50, 48, -9, 11, 41, 91, 141, 52, -20, 30, -10, 31, 21, 12, 19, 20, 42, 49, 19, 10, 1, -14, -14, -26, -52, -53, -28, 63, 71, 17, 48, 17, 28, 114, 168, 81, 33, 42, 27, -10, 18, 43, 39, 37, -26, -16, -21, -18, -17, -46, -6, 10, -2, -17, 12, 60, 58, 46, 70, -6, 18, 87, 157, 100, 87, 42, 41, 43, 42, 71, 57, 51, 16, -13, -6, 13, -26, -24, 0, -6, 6, 7, 54, 20, 51, -1, 7, -23, 20, 97, 103, 85, 93, 74, 19, 37, 78, 71, 33, 13, -30, -18, -8, -47, -46, -16, -15, -31, 16, -14, 22, -28, 21, 0, 51, -18, 18, 68, 91, 141, 125, 41, 31, 48, 36, 9, 3, -34, -26, -63, -61, -32, -24, -4, -8, -16, -8, 26, 23, -21, 34, -10, -1, -13, -36, 23, 89, 109, 119, 115, 58, 39, 8, -23, -15, -7, -10, -11, -36, -8, -14, -28, -38, -5, 30, 1, -13, -32, 18, -14, -15, -20, -45, 38, 98, 131, 88, 63, 94, 26, 16, -1, -14, 2, 17, -21, -2, -5, -9, -11, -67, -53, -29, -43, -30, 10, 21, 39, -2, 10, -10, 27, 20, 44, 11, 26, 35, 53, -16, 28, -6, 2, 2, -31, -48, -16, -24, -68, -90, -97, -88, -68, -47, 30, -37, 34, -12, -2, 14, 20, -39, -76, -64, -66, -53, -46, -44, -28, -60, -70, -113, -117, -84, -124, -153, -143, -102, -80, -84, -58, -34, -22, -10, -7, 14, -9, -10, -18, -8, 4, -54, -50, -37, -70, -43, -87, -67, -89, -26, 16, -73, -71, -58, -56, -30, -14, -23, -40, -3, 16, 6, 10, -10, -12, 9, 10, 19, -5, 9, 18, 12, 18, -12, -6, 21, 4, 12, -20, -32, -18, 1, -14, -9, 10, -16, 12, -17, -19, 2, -15, -4, 3, -1211, -11, 20, 6, 14, 16, 39, 15, 43, 45, 69, 107, 13, 5, 68, 63, 41, 23, 51, 42, 26, 28, 20, 32, 7, -18, 7, -20, 17, -1, -8, 2, 18, 22, 96, 80, 107, 121, 97, 62, 57, 90, 155, 83, 32, 67, 118, 127, 103, 89, 17, 1, -24, 29, -18, -15, -9, 15, 6, 25, 27, 25, 49, 70, 47, 77, 39, 36, 44, 32, 12, 10, 24, 53, 31, 21, 47, 44, 0, 31, 9, 43, -1, -1, -12, 20, 5, 0, 15, 40, -7, -23, 16, -2, -30, -15, -22, -14, -59, -47, -43, -48, -30, -27, -22, -39, -1, 60, 45, -16, -5, 21, -16, 8, -33, 2, 66, 32, 7, -42, -48, -60, -113, -68, -90, -70, -58, -80, -71, -69, -74, -80, -66, -14, -57, 3, -24, -102, -46, 6, 4, 20, -21, -11, 29, -6, -56, -94, -70, -114, -88, -54, -18, -36, -35, -49, -36, -73, -58, -56, -67, -46, -86, -60, -23, -111, -41, -17, 2, 4, -2, -12, 17, -55, -85, -95, -82, -97, -64, -31, -19, -25, -10, 25, 31, -31, -83, -94, -89, -108, -106, -51, -46, -105, -34, -25, 1, -19, -54, 11, 19, -23, -75, -96, -91, -24, -49, -40, -19, 1, 27, 60, 55, 18, -17, -98, -129, -177, -181, -145, -51, -75, 30, 14, -1, -26, -35, -51, -75, -30, -41, -34, -10, 16, -26, 22, -31, -9, 0, 6, 45, 39, 44, -8, -74, -157, -173, -109, -55, -57, 29, 27, -9, -25, 25, 36, -56, -41, 9, -11, -3, 41, 18, 19, -4, 15, -19, 6, 10, 36, 78, -8, -50, -74, -120, -77, -30, -92, -19, 1, 30, 18, -4, 44, 11, -18, 7, 37, 26, 2, 12, 12, -12, -30, -30, -39, 1, 41, 39, 40, -23, -55, -76, -14, -27, -57, -39, -35, 20, 15, -15, -70, -24, -13, 20, 45, 31, 27, 24, 5, -15, -16, -43, -59, -25, 47, 47, 9, -24, -40, -3, 4, 5, -58, -23, -2, 10, -41, -106, -21, -9, 26, 31, 46, 54, 44, 36, 5, -20, -3, -33, -15, -13, 32, 35, -16, -71, -69, -2, 8, -26, -5, -71, -14, -17, -8, -26, -9, 12, 53, 6, 40, 51, 18, 8, -9, -22, -8, -37, -3, -21, 44, 23, -24, -70, -36, -16, 4, 19, 29, 41, 20, -23, -24, -40, -27, -7, 0, 32, 5, 24, 3, 7, 17, 24, 18, 10, -15, -52, -20, -17, -54, -51, -50, 11, 24, 73, 50, 53, 10, 1, 10, -12, -72, -58, 35, 9, 3, 13, 18, 49, 40, 65, 48, 34, -2, -28, 10, -30, -45, 0, -13, 18, 35, 41, 34, 66, 37, 21, 15, -114, -121, -89, -23, 22, 31, 55, 30, 55, 27, 31, 28, 61, 102, 51, 43, 3, -9, -6, 25, 12, 22, 56, 47, 86, 52, 24, -4, -45, -63, -91, -63, -17, 19, 12, 31, -13, -22, -9, -12, 61, 69, 11, 32, -20, 4, 11, 19, 35, 35, 22, -28, 56, 68, 19, 40, -63, -140, -101, -116, -54, -23, -37, -3, -6, -30, -66, 22, 44, 34, 41, 29, 28, 9, 47, 25, 58, 34, -2, -26, -7, 66, 39, -47, -84, -172, -135, -97, -87, -61, -35, -29, -21, -13, 5, 22, 43, 39, 49, 10, 7, 30, 70, 35, 26, 21, 12, -10, -2, 59, -39, -40, -74, -97, -138, -153, -123, -72, -38, -8, 2, 48, 42, 35, 68, 39, -7, -5, 18, 26, 24, 32, 26, -33, -2, 29, 48, -1, 4, -26, -43, -103, -174, -207, -137, -54, -50, -44, -2, 34, 18, -17, -43, -29, -62, -38, -34, 5, 27, 25, 26, 17, 24, 21, 19, -32, -7, -4, -37, -90, -151, -204, -159, -106, -51, -35, -77, -119, -183, -148, -190, -136, -132, -113, -63, -42, -16, -51, 27, 24, 38, -61, -8, -3, 19, 19, -15, -49, -97, -125, -123, -40, 10, -3, 3, -13, -31, -62, -92, -85, -84, -49, -46, -36, -57, -28, 19, -16, 33, 19, -47, -18, 4, 6, -18, 10, 26, 24, 0, 61, 89, 97, 83, 63, 64, 79, 48, 49, 37, 74, 44, 80, 60, 76, 79, 63, 10, 40, -38, 6, -10, -4, 4, 17, 61, 54, 41, 89, 99, 102, 77, 25, 7, 19, 52, 5, 68, 145, 103, 74, 71, 98, 63, 39, 46, 39, -8, 8, -21, 19, -3, -5, -9, 54, 36, 63, 84, 66, 68, 93, 40, 7, 11, 90, 131, 63, 83, 66, 26, 64, 31, 10, 9, -10, 2, 4, -4, 17, -13, -5, -19, 5, -3, -7, 8, -6, 15, -2, 1, -6, -9, 16, 2, -2, -7, 11, 8, 17, 5, 18, 9, -7, 4, -4, -16, -1538, -6, 5, 12, -21, 37, 52, 50, 52, 68, 23, 38, 41, 51, 107, 25, 24, 0, 23, 38, 45, 39, 30, -12, -19, -1, 18, 18, 4, -19, 19, -2, 6, 50, 39, 49, 92, 56, 60, 26, 36, 10, 27, -12, 0, -10, 17, -33, 21, -21, -19, 2, -2, 17, 9, -5, 18, -11, 5, 45, -18, -29, -14, 27, 52, 64, 31, 37, 23, -22, -35, -36, -37, -138, -172, -146, -65, -60, -34, -2, 6, -10, -2, 21, -16, 11, 53, 74, 34, 26, 55, 58, 46, 38, 58, 15, -14, -10, -44, -95, -107, -90, -97, -86, -83, -70, -64, -22, -32, -77, -32, -3, -12, -18, 2, -14, 19, 55, 73, 56, 63, 71, 30, 24, 7, -20, -25, -32, -31, -55, -43, 16, -5, 13, 30, 58, -2, -58, -31, -18, 1, -22, -47, -23, 41, 27, 51, 61, 68, 47, 26, -11, 4, -41, -41, -36, -70, -42, -13, 1, 25, 12, 52, 107, 64, 43, -3, -8, -15, -11, -24, 0, 42, 30, 22, 72, 46, 57, 32, -7, 5, -17, -26, -49, -60, -28, -10, 17, -6, 13, 10, 50, 70, 36, 34, -4, 6, 7, 34, 48, 51, 20, 46, 13, 3, 28, -4, -20, 1, 7, -35, -13, -18, -17, -1, 13, 33, 33, 28, 24, 44, 54, -9, -47, 17, 18, 58, 44, 31, 37, 51, -18, -9, 15, -8, -33, -11, 15, 19, -1, -9, 10, 34, 6, 35, 55, -3, -17, 37, 34, -62, -10, -11, 51, -3, 62, 23, 20, 37, -29, -45, -20, -38, -9, -25, 49, 37, -4, -2, 18, 30, -3, -1, 17, -4, 15, 21, 62, -31, -30, 38, 50, 69, 54, -2, 5, -15, -45, -58, -84, -74, -17, -6, 19, 73, 62, 63, 44, 22, -3, -2, -8, 4, -2, 0, 8, -16, -49, 11, 54, 75, 15, 22, 0, 13, -42, -99, -85, -68, -11, -14, 9, 27, 48, 32, 18, -5, -33, -51, 15, 3, -15, -41, -31, -20, -48, -5, 41, 47, 19, -40, -73, -68, -71, -93, -82, -45, 26, -2, -11, 10, 37, -17, -23, -74, -43, -34, -40, -31, -97, -61, -27, -21, -22, -10, 34, 95, 20, -43, -65, -67, -92, -86, -20, 36, 7, 3, -34, 13, 20, -53, -79, -105, -110, -78, -55, -58, -134, -63, -58, 4, -35, -25, 50, 83, 51, -22, -63, -91, -97, -38, -1, 36, 30, 15, -26, 13, 2, -71, -75, -115, -102, -65, -44, -90, -92, -53, -45, 43, -5, 22, 32, 36, 53, 30, -110, -107, -52, 2, 42, 35, 26, 7, 8, -18, -122, -107, -124, -98, -54, -26, -60, -46, -6, -25, -50, 24, -9, -13, 45, 18, 3, -10, -87, -70, -40, 23, 60, 46, 29, -12, -23, -54, -82, -83, -7, -23, -26, -2, -17, 9, 25, -20, -96, -48, -34, -15, 53, 28, -21, -69, -71, -56, -46, -42, -4, 27, -4, -7, -63, -60, -34, -15, 30, 31, 43, 8, -32, 36, 2, -47, -43, -16, -56, 19, 3, 17, -26, -79, -26, -43, -86, -34, -5, -15, -33, -58, -16, 3, 46, 72, 51, 82, 30, -5, -29, -17, -24, -13, -7, -19, -23, 21, 8, 1, -82, -78, -44, -7, -71, -61, -43, -53, -42, -40, -17, 77, 86, 56, 41, 57, -9, -16, -22, -33, -1, 37, -24, -17, 62, -29, 34, -17, -83, -54, -37, -18, -8, -37, -97, -42, -58, 0, 24, 93, 93, 42, 55, 46, 5, -8, -4, 20, -29, 26, 0, 26, 42, 2, 1, -17, -55, -55, -17, -14, -24, -64, -45, 0, 0, 41, 49, 68, 49, 49, 63, 66, 32, -23, 21, 46, -8, 23, 13, 20, -17, -20, -18, -26, -7, -43, 5, 10, 23, 12, -8, -11, -15, -15, -30, -5, -7, 16, 18, 3, -11, 13, 7, 32, 12, 44, 23, 19, 4, -1, -15, -10, -26, -52, -27, -43, 1, 9, -24, -46, -78, -75, -81, -54, -22, -36, -30, 2, -4, 55, 21, 31, -24, 0, -9, 17, 10, -16, 18, -27, 18, 6, -36, -32, -67, -32, -51, -47, -80, -103, -104, -122, -53, -41, -38, -4, 20, -21, -33, -6, -20, -41, 28, 15, 16, 16, 8, 13, 37, 11, 15, -17, -46, -57, -99, -27, -46, -17, -53, -39, -47, -38, -21, -4, 37, -1, -20, -29, -6, -9, -3, 9, 6, -14, -10, -14, 13, 7, -12, -25, -35, -42, -21, -23, 30, 34, -7, -13, -26, -61, -39, -49, -36, -29, -13, -16, 2, -23, 13, 4, -13, 2, -15, -11, 17, 19, 19, 11, -17, -1, 10, 7, -12, 16, -2, 13, 6, 15, -18, -19, -11, 11, 6, 7, -2, 10, -16, -21, -7, 2, 157, -18, 1, 0, -9, 32, 26, 5, 30, 69, 65, 75, 76, 67, 91, 76, 42, 45, 49, 59, 22, 36, 47, 1, 19, 16, 14, 1, 14, 7, 19, -11, -1, 14, 63, 56, 124, 84, 113, 85, 103, 59, 163, 128, 120, 92, 70, 75, 50, 77, 53, 37, 29, -20, -3, 10, -20, -18, -31, -5, 40, 47, 37, 14, 19, 22, 1, 22, 22, 31, 57, 80, 97, 64, 125, 110, 98, 59, 70, 83, 23, 0, -8, -6, 12, 2, -16, -28, 19, 51, -1, -24, -13, -23, -31, 4, -17, 32, 81, 119, 113, 68, 149, 95, 97, 41, 53, 54, 41, 45, 19, 8, 10, 4, 32, 63, 66, 28, -3, -34, -14, -47, -15, 34, 36, 25, 32, 50, 68, 64, 71, 68, 88, 69, 78, 86, 18, 9, -43, 10, 19, -1, 0, 46, 62, 53, -18, -2, 11, -12, 17, 20, -2, 0, 21, 31, 19, 4, -6, 46, 40, 103, 118, 62, 31, -25, -30, -5, -19, -8, -34, 51, 85, 52, 35, 23, 36, 33, 17, -31, -10, -1, 1, 22, -8, 15, 15, 14, 16, 72, 48, 33, 8, -11, -7, -23, 2, 18, -23, 53, 68, 85, 78, 3, 35, 50, 2, -29, -33, -13, 8, 16, 46, 32, -4, 6, 30, 27, 67, 28, -14, -24, 26, 45, -20, -26, 16, 69, 44, 46, 20, 15, 36, 51, -16, -27, -41, -26, 15, 53, 11, -8, 29, -29, 21, 14, 52, -1, -33, -37, 49, 26, 18, -29, 67, 32, 39, 9, -4, -21, -7, 25, -11, -24, -20, -18, 33, 10, -27, 42, 31, -15, -34, 14, 29, 37, -47, -46, -31, 7, 37, 35, 23, -1, 40, 0, -58, -102, -13, -24, -45, -19, -41, -18, 10, 13, 40, -1, -26, -34, -31, 5, 46, 69, 14, -26, -32, 31, 9, 27, -30, -51, -2, -38, -71, -104, -73, -59, -26, -50, -66, -61, -11, 11, -21, -18, -16, -37, -44, -44, -13, 9, 53, -9, -70, -11, -9, 2, -10, 4, 4, -3, -80, -49, -32, -38, -3, -51, -45, -19, -4, -41, -68, -73, -23, -15, -26, -43, -29, -11, -15, -45, -69, -11, 1, 29, 24, -2, 21, 6, -29, -10, 1, -5, -23, -32, -27, -5, 8, -9, -61, -61, -43, -54, -20, -13, -11, -61, -32, 5, 22, 16, 18, -7, 54, 73, 9, -27, -15, -33, 30, -3, 5, -23, -3, -29, 47, 10, -51, -65, -14, -18, -4, 3, -37, -27, 10, 52, 9, -1, -1, 18, 90, 79, 57, 52, 4, -6, 21, 24, 21, 36, -8, 14, 76, -3, -22, 0, -19, 16, 11, 18, 2, -11, 36, 33, 34, 19, 16, 31, 60, 136, 158, 103, 75, 54, 70, 28, 75, 43, 29, 35, 58, 62, 48, 74, 58, 6, 25, 44, 55, 1, 44, 7, 38, -22, -3, 56, 92, 95, 180, 161, 93, 71, 55, 71, 19, 30, 15, 6, 43, 61, 86, 96, 82, 43, -15, 20, 94, 34, -8, 30, 55, 19, 30, 32, 69, 121, 158, 137, 143, 86, 70, 50, 66, 10, -30, -3, 40, 51, 70, 91, 87, 46, -2, 36, 60, 29, 0, 9, 18, 56, 3, 26, 44, 110, 141, 117, 106, 55, 68, 61, 37, -4, -29, 4, 16, 51, 98, 65, 25, 13, 42, 35, 50, -25, -15, -1, 4, 38, -38, -12, 23, 50, 30, 35, 7, 45, 33, 42, 30, -12, -2, 12, 42, 87, 109, 95, 83, 38, 13, 27, 13, -67, -46, 17, 37, -17, -8, 10, 6, -6, 7, -27, -15, 53, 41, 36, 50, 30, 53, 29, 70, 100, 140, 117, 59, -5, -14, 2, -22, -23, -82, -1, 4, -23, -14, -20, 19, 12, -46, -39, 20, -16, 21, -4, -28, -6, -18, -4, 10, 60, 74, 82, 12, -27, -53, -24, -61, -27, -78, 43, 30, -6, 20, -7, 39, 14, 7, -28, -30, -49, -77, -32, -11, -48, -20, 14, 1, -11, 17, 4, -67, -74, -51, -84, -47, -44, -25, 87, 30, 20, -3, -7, -27, 14, -42, -42, -28, -39, -35, 4, -3, -12, -4, -24, -38, -20, -7, -91, -86, -99, -74, -51, -60, -30, -8, 29, 33, -8, -15, -10, 6, 1, -31, -40, -56, -33, -31, -22, 15, 9, -23, -38, -101, -92, -59, -91, -43, -26, -37, -12, -73, -23, 1, 25, 17, -9, 20, -1, 16, 0, 15, -49, -59, -63, -48, -63, -57, 35, 40, 59, 13, 15, 13, 3, -27, -25, -8, -15, 1, 0, -8, -15, 3, 11, -13, -7, -8, -13, -3, 15, -2, -19, -16, -19, -6, -11, -13, -12, -4, 7, -19, -8, -21, -7, -5, -21, -12, 17, -8, -5, 1, 5, -11, -1359, 17, -14, -13, 4, 26, 31, 50, 63, 54, 59, 50, 78, 83, 89, 56, 43, -2, 37, 34, 29, 37, 13, 9, 8, -8, -3, 12, 7, 6, 10, 12, 34, 50, 22, 30, 20, 16, 16, 19, 24, 35, 85, 1, 11, -13, 12, 27, 81, 107, 50, 44, 26, 19, 16, -7, -17, -13, 31, 54, -36, -69, -21, -6, 50, 13, 0, -22, -28, 3, 38, -2, -35, -68, -75, -1, 23, 6, 10, 62, 18, -36, 8, -15, -8, -7, 55, 44, 15, 47, 32, 116, 72, 69, 39, 19, -1, -12, -42, -79, -80, -61, -20, -30, -43, -51, -36, 10, 56, -35, 5, -1, -3, -10, -2, -24, 33, 26, 34, 68, 78, 34, 53, 16, -18, -41, -64, -40, -11, -11, 0, -28, -34, -16, -13, -5, -13, 2, -18, 20, 6, 11, -38, 2, -1, -15, 19, 43, 32, 3, 18, -2, -22, -62, -57, -60, -39, -29, -2, -16, -14, 9, 10, 27, 14, 88, 59, -19, 17, 17, -29, -17, 0, 10, 12, 16, 20, 5, 8, 8, -15, -51, -44, -54, -42, -33, 14, -20, -11, -26, -32, 18, 19, 48, 71, 42, -1, -4, 53, 12, 12, 5, -9, 25, 41, 27, -8, 3, 4, -31, -17, -10, -33, -16, -21, -9, 5, -9, -25, -31, 55, 40, 13, -25, -19, 10, 57, 31, -66, -7, 6, 24, 28, 13, -6, -9, 11, 27, 15, 25, -70, -75, -51, -40, -31, -12, -41, 9, 45, 21, -9, -18, 5, 18, 7, 20, 0, 11, 16, 6, -6, 21, 29, 2, 12, 10, 19, -1, -50, -65, -80, -68, -63, -42, -19, -13, 29, 56, 8, -4, 27, 11, 68, 62, -21, -9, -11, 31, -17, -14, 8, 34, 15, 42, 61, 84, -3, -59, -61, -92, -49, -40, -13, -30, 26, 16, 4, -19, 18, 48, 110, 26, 13, 2, 4, 26, -11, -31, -3, 38, 67, 85, 74, 54, 19, -29, -49, -30, -34, -10, 1, -26, 1, 14, 12, -15, 15, 59, 43, 7, -34, -25, -51, -52, -38, -3, 35, 76, 83, 90, 60, 47, -5, -71, -55, -71, -31, -48, -46, -14, 44, 48, -2, -4, -1, 45, 109, 95, -14, -38, -52, -82, -47, 27, 37, 37, 40, 15, 32, 11, -37, -19, -48, -36, -39, -37, -35, -48, 56, 66, 28, -19, -39, 46, 99, 105, 35, -83, -120, -86, -47, -3, 14, 27, 13, 30, 49, -13, -30, -6, 18, 13, 29, -32, -28, -28, -6, 58, 18, -13, -8, 72, 61, 51, -35, -126, -150, -72, 16, 38, 41, 9, 22, 35, 34, -47, -28, 14, 26, 0, -15, -30, -53, -10, 25, 49, 35, 14, -13, 37, 27, -52, -165, -175, -121, -60, 54, 92, 64, 19, 45, 36, -13, -39, -8, -8, 1, -19, -15, 4, -5, 50, -1, 112, 60, -22, 5, 41, -11, -57, -194, -175, -120, -26, 10, 71, 74, 52, 55, 35, -8, -18, -30, -20, -19, -11, 4, 35, 29, 69, 32, 124, 67, 18, -24, 1, -48, -103, -188, -145, -101, -30, 18, 58, 71, 43, 70, 67, 5, 16, -42, -51, -3, -23, -5, 24, 52, 48, 29, 86, 48, 16, -11, -3, -47, -121, -180, -175, -88, -29, 13, 46, 38, 20, 22, 13, 2, 19, -38, -56, 3, -2, -12, 36, 16, 9, 73, 75, 19, 44, -42, -15, -15, -44, -105, -125, -64, -32, 18, 24, -15, 25, 21, -6, -19, 23, 4, -25, -20, -21, 2, -1, -2, -40, 71, 60, 14, 11, 2, -16, -19, -60, -111, -111, -94, -13, -22, -4, 8, 32, 43, -18, 26, 28, 22, -17, 18, 28, -7, -2, -9, -11, 6, 70, 3, 4, 15, -48, -59, -60, -90, -63, -29, -45, -65, -29, 13, -11, 10, 18, -6, 34, 5, -2, -16, 3, -17, 0, 0, 31, 28, 23, 18, 17, 17, -41, -76, -82, -73, -126, -40, -76, -80, -44, -16, -8, 11, 8, 1, -1, -14, -8, -39, -37, -5, -12, -8, 16, -42, -8, 34, -10, 16, -15, -38, -10, -79, -34, -18, -74, -88, -50, -46, -10, -21, -3, -54, -31, -30, -26, -24, -12, -76, -53, -37, -8, -58, -43, 30, -5, 4, -10, 5, -3, -25, -69, -75, -88, -83, -108, -34, -37, 30, -34, -50, -32, -35, -30, -36, 11, -29, -53, -44, -25, -21, 4, -17, -5, 10, -8, -17, 7, -20, -26, -24, -47, -44, -29, -58, -57, -22, -12, -3, -87, -43, -58, -22, -54, -58, -35, -21, -15, -4, 20, -16, 13, 7, 5, -6, 12, 11, -11, -5, -10, -11, -8, 0, -19, -1, -12, 1, -7, -25, -10, -11, -18, 16, 8, 3, -19, 4, 11, 20, -9, 9, 967, 12, -8, 0, -1, -11, -65, -30, -36, -53, -78, -69, -72, -53, -122, -48, -62, -33, -62, -38, -55, -56, -41, 14, 2, 2, -4, 17, 15, -8, 13, -5, -25, -11, -85, -98, -127, -100, -94, -79, -101, -102, -154, -112, -58, -62, -128, -134, -128, -95, -86, -45, 6, 13, 19, 20, 19, -13, 16, 2, -9, -25, -11, 1, -44, -77, -36, -56, -54, -26, -40, -39, -44, 1, -5, -45, -94, -71, -69, -54, -34, 24, -1, -5, 9, 4, -8, -14, -39, -23, -6, 22, 3, 11, 22, -9, 28, 16, 25, 17, 45, 59, 34, 55, 27, 12, -30, -75, -86, 19, -5, -19, -20, -19, 35, 3, -52, -22, 25, 84, 81, 74, 47, 27, 43, 52, 54, 69, 74, 99, 89, 116, 90, 74, 29, -33, -33, 46, 32, -11, -9, -5, 23, -18, -25, 19, 48, 91, 38, 88, 41, 54, 7, 26, 36, 51, 50, 113, 71, 88, 78, 100, 79, 8, -19, 14, -16, 6, -3, -6, 27, -8, -38, 14, 49, 53, 46, 42, 33, 15, -8, -3, 24, 13, 45, 67, 24, 93, 86, 112, 93, 18, -2, 5, -26, -15, 2, -14, -20, -31, -8, -30, 20, 33, -3, -12, -17, -8, -11, 2, 12, 20, 30, 5, 9, 56, 66, 86, 118, 36, -12, 12, 46, 19, -12, -11, -29, -53, 47, 9, -10, -16, -1, -71, -38, -8, -28, 19, 8, 34, -31, -13, -40, 9, 24, 65, 104, 32, -2, 4, 14, -3, 11, 2, -75, -101, 64, 10, -47, 0, -2, -39, -34, -2, 29, 23, 49, 56, -12, -15, -63, 14, 0, 29, 51, 7, 12, -27, -34, 7, -19, -38, -75, -70, -7, 29, -36, -19, -28, -48, -13, 26, 69, 57, 33, -1, -38, -32, -12, -2, 32, 17, 19, 1, 6, 1, 3, -28, -8, -16, -62, -15, 2, -9, -42, -33, -34, -56, -10, 37, 37, 47, 53, 39, 31, 3, -17, 5, 43, 23, 20, 2, -15, 7, -5, -1, -27, -22, -16, -23, -24, -6, -22, -62, -57, -57, -30, 20, 41, 11, 7, 25, 30, -20, -19, 22, 46, 46, 34, 2, 15, -5, 51, 12, 11, -14, -78, -55, -52, -82, -32, -43, -47, -34, 13, 15, 14, 11, 4, -1, 10, 29, 21, 29, 27, 40, 8, 8, -31, -52, -58, -19, 13, 0, -45, -44, -51, -43, -27, -19, -21, 10, -6, -43, -52, -17, -41, 30, 57, 59, 46, 42, 24, 17, -29, -9, -52, -47, -45, -4, 4, -49, 1, -21, 3, -58, -45, -9, -13, -24, -61, -73, -58, -32, -22, 54, 43, 36, 49, 18, 6, -22, -24, -32, -84, -62, -40, -30, 11, -7, 78, 93, 29, -49, -45, -13, -39, -19, -57, -57, -25, 15, -25, -51, -20, -5, 31, -8, -3, -48, -18, -62, -53, -21, -75, -16, 0, -5, -13, 89, 80, 13, 0, 22, 15, 19, -35, -16, -2, 9, -38, -86, -15, -6, -5, -8, -25, -39, -62, -22, -18, -13, -32, -40, -27, -26, -11, 94, 94, 101, 40, 75, 66, 53, 4, -19, 20, -8, -61, -37, -39, -50, -48, -23, -27, -15, 10, -28, -32, -21, -2, -57, -11, 7, 50, 120, 112, 121, 130, 127, 94, 90, 68, 43, 54, 16, -34, -56, -37, -27, -58, 5, 1, -3, 21, 34, -27, -7, 0, -23, 21, 22, 41, 82, 132, 167, 198, 159, 153, 136, 151, 95, 6, -12, -82, -65, -54, -7, -47, -20, -18, 18, -1, 61, -28, -29, -65, -23, 15, -3, 37, 44, 127, 190, 193, 166, 170, 179, 135, 89, 44, 25, -33, -32, -32, -50, -23, -10, 34, -3, 12, 31, -58, -45, -37, 9, -1, -12, 8, 17, 83, 120, 153, 137, 150, 99, 167, 196, 177, 139, 133, 83, 48, 22, 28, 7, -6, -27, -27, -78, -87, -58, -1, -6, -8, -18, -6, 12, 58, 82, 97, 34, 64, 53, 42, 94, 111, 106, 87, 70, 49, 21, 3, -48, -47, -42, -81, -54, -64, -55, 21, 14, -14, -11, 10, -23, -9, 3, 5, -33, -33, -27, -71, -23, -23, -46, -37, -68, -79, -91, -71, -99, -119, -69, -78, -46, -43, -51, 4, 1, -11, -4, 7, -34, -30, -47, -46, -74, -61, -68, -63, -53, -45, -58, -49, -29, -75, -159, -139, -118, -89, -52, -38, -15, -30, -4, -11, -9, 2, -1, 7, -13, 13, -44, -61, -52, -62, -46, -89, -62, -43, -26, 1, -4, -41, -52, -34, -43, -38, -52, -42, 3, -23, -2, -15, -7, -8, 13, 16, -4, 20, 11, 6, -5, -15, 5, 8, 9, 2, -9, -17, 6, 11, -12, 13, 16, -1, 21, -13, 8, -21, 7, -1, 12, 16, 608, 5, 9, -11, -16, 36, -46, -31, -48, -51, -42, -61, -65, -80, -94, -7, 5, -31, -35, -19, 16, 1, -10, 19, -19, 5, 9, -3, -1, 11, 1, -8, -46, -54, -50, -47, -62, -32, 1, -25, -26, -51, -66, -19, 21, -13, -41, -78, -41, -67, -87, -93, -61, -1, -10, -14, 7, -7, -30, -11, 48, 27, -7, -66, -52, 26, 33, 67, 57, 25, -30, 14, 21, 31, 35, 46, 31, 21, 15, -24, -40, -36, 7, 2, -5, 16, -14, -59, -39, -48, -50, -19, 14, 55, 70, 42, 76, 91, 66, 66, 23, 12, -4, 19, -9, -7, -9, 10, 52, 76, 46, 2, 14, 2, 24, -53, -83, -65, -21, 10, 31, 57, 81, 60, 74, 50, 63, 75, 26, 30, 13, -19, -40, -53, -16, 30, 52, 99, 83, 19, -12, -21, -10, -91, -103, -2, -21, 17, 69, 87, 65, 63, 69, 45, 48, 43, 10, 19, -9, -14, -57, -36, -45, -36, -8, -8, -15, 10, 14, -16, -43, -118, -88, -19, -13, 43, 62, 74, 82, 29, -2, 35, 77, 33, 42, 3, -20, -12, -14, 21, -9, -65, -53, 17, -1, 7, 0, -10, -89, -85, -69, -5, 36, 23, 60, 0, 17, -14, -31, 23, 23, 4, -7, -40, -33, 6, -15, -18, -2, -19, -34, -1, -36, 34, -10, -39, -89, -60, 10, 21, -13, -1, 8, -13, -18, -48, -41, -24, -6, 25, 26, -29, -9, -38, -32, -53, -56, -20, -16, -5, 8, 24, 7, -51, -51, -59, 10, 3, -41, -47, -20, -37, -54, -71, -51, -52, -9, 38, 46, 44, 21, -7, -27, -43, -10, -29, -43, 38, 24, 30, -25, -91, -132, -59, 4, 6, -74, -72, -35, -14, -36, -64, -82, -77, -16, 45, 80, 24, -27, -31, -34, -61, -23, 8, 34, 50, 19, 42, -10, -74, -176, -46, 1, -8, -73, -71, -40, -23, -51, -95, -79, -58, 48, 95, 50, -5, -21, -28, -69, -85, -44, -12, 28, 38, 43, 50, -29, -44, -101, -23, -43, -64, -115, -53, -65, -23, -53, -92, -50, 15, 58, 46, 9, -14, -24, -41, -75, -42, -29, -18, -2, -30, 94, 35, 22, -47, -96, -102, -60, -117, -160, -88, -65, -17, -22, -42, -11, 46, 66, 27, 22, -14, -24, -38, -62, -61, -44, -49, -18, -6, 39, 35, 7, -29, -61, -52, -106, -146, -145, -58, -19, -7, -35, -60, -3, 73, 62, 52, 38, -13, -38, -33, -49, -56, -21, -35, -12, 26, -14, 9, -18, -35, 21, 0, -89, -98, -108, -35, 4, -8, -44, -11, 60, 140, 115, 43, 12, -19, -15, -8, -23, -8, -35, 20, 29, 35, -32, -11, -28, 34, 112, 56, 26, -3, -43, -36, -15, -35, -28, -18, 64, 142, 135, 64, 23, -9, -35, -48, -9, -17, -17, -18, 53, 36, -37, -33, -22, 49, 84, 82, 67, 8, -30, -5, 1, -35, -42, -23, 41, 114, 82, 32, 0, -26, 3, -7, 10, 29, -7, -26, 28, 28, -47, -67, -3, -5, 87, 116, 32, -1, 14, -1, -41, -5, -15, -11, 25, 63, 38, 19, 28, -5, -53, -9, 26, 27, -12, -28, -2, 2, 28, -50, 17, 9, 21, 38, 14, 1, 16, 7, -13, -5, 12, 14, 1, 13, 21, 22, -2, 1, -44, -23, 2, 34, 5, 31, 7, 46, -48, -57, -16, 24, 27, 46, 11, 20, -3, -36, 3, -8, -17, -7, -17, 20, 22, -8, -14, -44, -12, 14, 15, 6, -48, -5, 31, 26, -63, 50, -12, 16, 72, 124, 107, 50, 27, 11, 14, 25, -16, -6, -17, -1, -16, 12, 6, -22, 10, 12, 15, -8, 5, -3, 9, 19, -5, 19, 3, 12, 77, 44, 39, 60, 45, 55, 62, 43, 31, 22, 50, -4, 11, 0, 7, -31, -10, 28, -4, 16, -5, -17, -6, 29, -25, 18, 14, 17, 52, -7, 32, 44, -14, 58, 29, 43, 33, 38, 30, 56, 41, 16, -14, -9, 11, 23, 0, 2, -33, 30, 21, 33, 12, 8, 12, -8, -3, -35, -8, -17, -3, 18, 43, 12, 43, 22, 33, 28, 30, 33, 1, -4, 4, 9, 53, 24, 11, 36, 21, 44, 11, 4, -15, -8, -8, -15, -35, -22, -1, -50, -13, 14, 46, 37, 47, -2, 1, 1, -19, -5, -8, -51, -14, -12, 17, -8, 14, -15, 13, -19, 10, 15, 18, 2, 0, 37, 47, 64, 77, 40, 73, -30, -22, 20, 4, 40, 41, 61, 20, 36, -4, 47, 35, 7, -11, 13, 7, -16, -8, -16, 3, 20, -18, 11, 6, 15, 0, 1, -18, -16, 1, 13, -18, -9, -3, -3, -10, -18, 6, 15, -2, -17, 10, -9, 2, -3, -16, -92, -2, 17, 9, -17, -19, 18, 16, -15, 16, 22, -21, -23, 31, 36, -70, -16, -15, -16, -22, -14, -13, 6, -36, -25, -19, -12, -7, -18, 19, 0, 5, 4, 33, 48, 66, 72, 15, 7, 27, 19, 46, 67, -10, 5, 15, 5, -19, 34, 62, 96, 76, 74, -14, -3, -13, 12, -1, -24, 29, -38, -26, 32, 49, 56, -13, -4, -16, -30, -15, 4, -42, -48, -44, -47, -50, -81, -97, -10, 38, -41, -20, 11, -2, -9, 8, 9, 11, 10, 38, 65, 103, 79, 4, 5, 38, -3, 23, -15, -3, -12, -35, -36, -29, -33, -18, -25, -25, -60, -108, -70, 15, -14, -6, -52, -3, 59, 2, 55, 57, 42, -1, 27, 44, 15, 11, 4, -12, -10, -18, -33, -33, -21, -6, 6, -15, -85, -60, -72, -9, 19, -8, -24, -6, 53, 0, 26, 36, -7, -30, 4, -15, 5, -11, -14, 8, 13, -22, -32, -42, -10, -47, 6, 23, -35, -28, 14, 13, -12, -5, 47, 16, 48, 8, 17, -7, 4, -25, 4, -6, 40, 13, -5, -22, -16, -39, -34, -67, -47, -54, -4, 21, -19, -27, 5, 4, 9, -11, 66, 35, -1, -22, -18, -28, -10, 0, -11, 2, 17, 33, 25, -1, -21, -39, -47, -59, -49, -49, -36, -2, 24, -33, 28, 24, 4, 12, 83, -10, -10, -40, 16, 13, 17, -3, -8, 35, 39, 53, 0, -86, -66, -6, -27, -27, -27, -3, -24, -31, -28, -32, -27, -19, 6, 43, 7, -5, -42, -66, -4, -7, -2, -9, 13, 47, 75, 65, -17, -130, -108, 1, 11, -32, -19, -21, -12, -13, 10, -69, -58, -7, -15, 20, 36, 1, -68, -66, 24, 26, 6, 17, 41, 63, 87, 15, -97, -129, -87, -39, -6, -37, -7, -14, 21, 52, 12, -74, 8, -34, 13, 66, 89, -3, -56, -26, 42, 7, 44, 6, 63, 109, 42, -22, -129, -121, -55, -6, -28, -15, 51, 85, 78, 111, 27, -51, -24, -35, 10, 46, 117, 0, 5, 16, 50, -2, 26, 24, 42, 97, 25, -106, -148, -61, 10, -16, -4, 39, 19, 83, 75, 138, 122, 24, -22, -23, -1, 55, 75, -7, 57, 39, 31, 11, 11, 28, 52, 37, -33, -103, -102, -37, -2, -13, 32, 35, 41, 117, 111, 139, 151, 41, -73, -8, -5, 32, -34, -33, 21, 48, 14, -13, -9, 21, 45, 38, -54, -98, -80, -42, 9, 24, 37, 37, 33, 67, 75, 73, 75, 9, -41, -3, 6, -42, -74, -97, -3, 18, 26, -9, 34, 20, 37, 8, -60, -78, -108, -63, -20, 6, 25, 20, 25, 1, 55, 19, 30, -22, -20, -6, -6, -44, -115, -108, -61, -1, 12, 37, 14, 14, -14, 4, -1, -53, -103, -73, -7, 10, 38, -22, -4, -20, 23, 34, -40, -52, -48, -2, -10, -19, -92, -71, -51, 17, -8, -6, 3, 3, 5, 47, 24, 1, -17, -6, -9, 3, -14, -39, -41, -22, 33, 36, -23, -31, -14, -16, -26, -9, -72, -170, -40, -16, -51, -14, 1, -6, 13, 38, 53, 38, -6, -1, -20, 6, -19, -41, -16, 18, 5, 31, -44, -64, -49, -17, -6, -8, -44, -105, 0, -30, -45, -2, -2, -20, 1, 32, 61, 74, 24, -19, -22, -34, -26, -26, -29, -41, 8, -12, -31, -67, -29, -46, 44, -20, -62, -76, -18, -11, 9, 8, -1, 14, -4, 24, 34, 39, 31, 41, 36, -8, -15, -37, -42, -17, 10, 6, -20, -27, 36, -85, 8, -27, -113, -147, -108, -60, 10, 10, 15, 10, 1, 9, -24, 2, 4, 38, -12, 3, -1, -58, -44, -16, 3, -18, -33, 7, -13, -47, -2, -29, -76, -90, -78, -75, -18, -7, -27, -24, 27, -10, -41, 29, -1, 27, -4, -2, -1, -46, -24, -30, -15, -55, -18, -3, -30, 3, 0, -28, -40, -81, -75, -18, 13, -3, -2, -12, -7, 11, -38, 3, 4, -11, -28, -23, -43, -20, -15, -5, -34, -60, -67, -30, 4, 7, -15, 11, -41, -22, -86, -82, -56, -31, -17, -7, -22, -9, -38, -25, -27, -26, -65, -57, -60, -44, -81, -30, -31, -44, -25, -1, -13, -17, -9, 16, -20, -26, -24, -49, -81, -59, -71, -113, -121, -127, -85, -127, -82, -79, -111, -161, -103, -91, -87, -67, -62, -12, -34, 20, -25, -8, 19, -13, 18, 16, -15, -26, -37, -48, -62, -62, -60, -15, 12, -1, -11, -34, -31, -47, -60, -78, -41, -67, -32, -28, -3, 2, -14, -7, 19, -17, 6, 4, 6, 21, -4, -14, 10, 19, 11, -13, -18, -2, 17, -13, -5, 1, 14, 20, 8, 7, 14, -9, 15, -2, 4, 12, 19, 779, 17, 14, 10, -2, -16, -7, -10, 4, 13, -14, -66, -15, 35, -5, -42, -5, -16, -26, -33, -75, -61, -46, -22, 6, -1, 4, 5, 2, -21, -20, 15, 3, -13, -50, -32, -6, -54, 33, 31, 3, -20, -1, -15, 9, -7, -26, 14, 39, 6, 4, 4, 47, -17, -5, -12, -11, 1, 12, -28, -46, -17, -69, -5, 13, 5, 31, 27, 40, 67, 34, -3, -68, -20, -20, -84, -92, -45, -17, -21, 8, 22, 8, -10, 2, -10, -48, 3, 2, 56, 30, 40, 100, 68, 15, -35, 20, 9, -20, 4, 1, -32, -68, -27, -44, -58, -58, -98, -78, -72, -12, 17, -4, -15, -49, 43, 19, 46, 52, 55, 36, -2, -29, -31, -23, -36, -1, -12, -48, -88, -65, -39, -26, -21, -50, -61, -43, -61, -41, 19, -4, 10, -14, 60, 66, 8, 47, 26, -40, -40, 0, -42, -9, -19, -14, -57, -67, -54, -47, -45, -29, -16, -14, -22, 22, -6, -39, -15, -16, 2, 17, 29, 16, 4, 15, -16, -26, -17, -6, 4, -45, -41, -59, -43, -64, -60, -19, -22, -48, -82, -83, -40, -16, -53, -45, 1, 7, -6, 23, 29, 26, -13, -32, -22, -15, -23, -28, -47, -41, -37, -49, -20, -28, -6, 0, 2, 14, -14, -81, -67, -75, -51, -24, -18, -5, 44, 36, -8, -27, 13, -2, -22, -19, -6, -26, -55, -65, -32, 8, 66, 63, 80, 86, 67, 91, 33, -3, -77, -52, -36, -37, -37, -3, 40, 12, 35, 10, 11, -46, -61, -30, -30, -44, -17, -22, 13, 56, 161, 172, 143, 141, 155, 129, 81, -14, -62, -87, -7, -23, -22, -35, -18, -28, 110, -3, -50, -70, -53, -46, -48, -44, 20, 64, 55, 119, 126, 134, 84, 139, 183, 162, 90, 37, -46, -108, -61, -10, -3, -17, 4, -32, 63, -27, -54, -101, -91, -59, -52, -27, 59, 63, 65, 32, 18, 31, 49, 91, 100, 119, 69, -4, -56, -89, -13, 8, -23, 18, 8, -32, 73, -72, -47, -39, -60, -79, -9, 0, 81, 65, 38, 20, 6, 1, 34, 25, 64, 57, 9, -27, -14, -76, 22, 37, -18, 11, 43, 34, 69, -63, -22, -37, -63, -70, -15, 33, 67, 58, 25, -2, 13, 25, 60, 5, -2, -10, -36, -31, 3, -42, 3, -14, -6, -16, 49, 29, 82, 15, 56, 16, -22, -53, -36, 28, 43, 62, 54, 0, 9, -3, 2, -13, 5, -13, -48, -44, 27, 5, -16, -7, 8, 14, -4, -26, 55, 94, 21, -14, -21, -52, -32, -23, 58, 63, 56, 14, 16, 27, -5, -19, 28, 19, -28, -26, 19, -17, -13, -18, 9, 15, -13, -60, -9, 45, 13, 6, 17, -27, -7, -9, 16, 73, 70, 47, 23, 27, 6, 26, 29, 0, -5, -18, 4, -16, -47, -67, 19, 20, -46, -84, -93, 4, 23, 12, -2, -16, 7, 15, 29, 50, 40, 34, -18, -5, 0, 5, 16, -15, -7, 21, 10, -7, -88, -40, 9, -21, -16, -5, -95, -35, 11, -3, -14, 14, -15, -23, -18, 7, 2, -21, -22, -14, 0, 12, 11, -29, -22, 32, 3, -29, 8, -7, 0, 3, 17, 14, -46, -13, -1, 12, -10, -48, -18, -32, -8, -21, -10, -38, -3, 4, 29, -12, 18, 7, 18, 15, -4, 37, -5, -2, -3, -13, -13, -35, -39, -15, 24, 24, 3, -30, -40, -8, -24, -10, 9, -48, -32, -33, 6, -17, 2, -3, -17, -13, -31, -17, -44, 6, -40, 7, -10, -31, -31, -34, -18, -19, -26, -45, -32, -29, -35, -19, -34, -17, -20, -1, 11, 12, 14, 5, -2, -43, -55, -4, -27, -25, -33, -6, 6, -30, -15, -23, -39, -12, -12, -25, -11, -45, 3, -10, -14, -16, -27, 9, 34, -8, -11, 14, -23, -44, -83, 6, -51, 19, 14, 12, 24, -40, -14, -23, 28, 4, 1, 24, -37, -42, 41, 29, -9, 23, -14, -6, -7, 3, -4, -28, -29, -15, -25, -24, -38, -38, -17, 3, 15, -15, 37, -8, 22, 67, 33, 0, 6, 1, -18, -25, -15, -20, -37, -41, 0, -6, -8, -37, -2, 0, 16, -12, -24, -3, 19, 4, -14, 12, -4, 32, 15, 11, -7, -10, -16, -19, -47, -50, -33, 16, 67, 61, 37, 26, 52, 38, 39, 54, -3, -16, -8, 8, -4, -17, 0, -11, -12, -16, -6, 9, -5, -7, 15, 11, 44, 51, 0, 21, 59, 33, 21, 35, 42, 43, 31, 34, -18, 17, 17, 4, -6, -9, 18, -16, -18, 10, 18, -16, 3, -14, -11, 7, 14, -14, -19, -4, -13, -4, 12, 6, 7, 12, 3, 19, -7, -16, -7, 18, -6, 9, -147, -12, 15, 1, 12, 32, 80, 89, 33, 45, 40, 39, 104, 113, 125, 69, 37, 17, 27, 60, 20, 26, 33, 16, 8, -10, 9, -11, -13, 16, 18, 19, 41, 39, 43, 47, 68, 21, 36, 15, 44, 77, 119, 48, 17, -15, 33, 65, 102, 110, 109, 104, 50, 14, -8, 10, 7, 8, 2, 1, -41, -33, -21, 28, 38, -8, 45, 30, 3, 18, 0, -46, -16, -5, -8, -9, 31, 21, 24, 62, 57, -10, 5, 3, -16, -3, -7, 23, 4, 21, 25, 62, 49, 40, 13, 35, 2, 7, -15, -45, -48, -2, -12, -38, 8, 21, 22, 23, 17, -84, -8, -3, -9, -15, -19, -7, 4, 44, 29, 27, 22, 19, -3, -24, -4, -5, 4, -4, 0, -15, -29, -18, 3, -31, -20, -53, -33, -101, -63, -18, -16, -19, -58, 8, 6, -17, -18, -36, -43, -34, -28, -41, -30, -37, -6, -31, 12, -6, 35, 26, 28, -40, -38, -88, -43, -87, -68, -10, 11, 3, -34, 3, 9, -27, -70, -60, -52, -5, -42, -27, -26, -34, -34, -10, -7, -18, 8, 48, 1, -91, -113, -34, -57, -136, -35, -36, -11, -13, -16, 31, 0, -69, -72, -74, -65, -36, -60, -60, -11, -54, -28, -24, -21, -18, -8, -46, -28, -104, -131, -84, -77, -128, -58, -31, 2, -40, -6, -16, -105, -128, -123, -77, -59, -15, -45, -55, -40, -36, -18, -33, -40, -19, -47, -78, -68, -80, -90, -72, -42, -46, -34, 7, -21, -7, 17, -41, -137, -159, -79, -56, -79, -57, -43, -41, -31, -37, 7, -67, -71, -53, -92, -112, -94, -70, -45, -48, -32, -44, -44, 5, 44, -59, -14, -4, -129, -114, -58, -68, -72, -70, -21, -16, -35, 15, -6, -57, -73, -102, -77, -82, -55, -9, -17, -4, -13, -62, -32, -3, -14, -52, -46, -89, -128, -70, -25, -40, -6, 6, 20, 33, 20, 4, -16, -68, -69, -68, -51, -88, -42, 23, 24, 3, 39, -37, -34, -37, 25, 3, -28, -50, -188, -48, 39, 37, 35, 57, 48, 72, 15, 4, -21, -56, -47, -15, -26, -82, -26, 10, 36, 35, 27, 54, -38, -11, -21, 12, -6, 9, -113, -25, 34, 93, 81, 85, 56, 25, 44, 46, 10, -27, -11, -32, -20, -16, 15, 68, 64, 54, 83, 37, 27, 15, -18, 18, 26, -38, -47, -59, 66, 74, 49, 35, -1, 28, 53, 61, 7, -56, -40, -2, -24, 5, 32, 70, 74, 70, 105, 21, 75, 40, -26, 50, -39, -55, -104, 1, 40, 57, 64, 25, 19, 12, 56, 72, -17, -82, -45, 35, 37, 24, 86, 58, 91, 48, 42, 13, 66, 47, 4, 38, -66, -48, -104, -57, 38, 26, 43, 11, 27, 51, 42, 49, -20, -33, 21, 41, 56, 61, 60, 58, 50, 59, -7, -3, 62, -16, 17, 15, -75, 8, -75, -34, -2, 27, 3, -15, 11, 17, 10, 25, -21, -34, 28, 48, 11, 33, -1, 18, 31, 55, -6, -3, 1, 37, 2, 36, -15, -31, -12, -23, -2, 9, -31, -18, 23, 9, -19, 20, 0, -34, 0, 6, 28, 3, 7, 10, 18, 11, -16, -8, 29, 37, -35, -17, 17, 35, 16, 17, -20, -19, -16, -28, -9, -16, -23, -6, -1, -41, -14, 0, 10, 7, 28, 8, 26, 16, 17, 24, 63, 42, -28, -34, 62, 22, 39, 13, 11, -18, -10, -6, 7, -1, 25, 16, 21, 41, 35, 4, 3, 46, 11, -19, 9, -13, -8, 73, 85, -48, 21, 5, -1, 1, 24, 5, -5, 7, -35, -23, 23, 44, 19, 14, 41, 7, 22, 43, 2, 26, 37, 5, -11, 0, 13, 26, -2, -23, 5, -27, -44, 12, 3, 1, -50, -58, -78, -74, -42, -67, -55, -37, -47, 17, -5, 6, -37, -21, -14, -73, -65, -38, -60, -8, -19, 9, 10, -24, -56, -19, 25, -5, -16, -40, -154, -195, -154, -183, -186, -237, -200, -130, -117, -123, -142, -157, -111, -100, -90, -55, -63, 8, 8, 1, 18, 5, 1, -31, -5, 18, -16, -69, -88, -74, -59, -121, -207, -195, -213, -178, -169, -129, -96, -74, -113, -138, -73, -49, -59, -20, 10, -17, 18, -5, -12, -26, -10, -34, -27, -22, -78, -113, -53, -81, -97, -111, -108, -144, -116, -85, -80, -62, -94, -76, -32, -23, -29, -19, -3, -2, -10, 0, -10, 11, -1, -47, -55, -33, -63, -21, -42, -74, -49, -42, -3, -53, -67, -45, -32, -55, -61, -20, -30, -12, 20, 21, 6, 5, -4, 6, -3, -6, 17, 0, -20, -5, 7, 12, 12, -15, -10, -18, 10, 11, -21, 11, 17, -4, -8, 19, -9, 7, -18, 15, -17, 5, 4, 2058, 11, 10, -11, 15, -32, -27, -5, 3, -45, -30, -26, -60, -37, -71, -47, -20, -40, -66, -37, -37, -27, -30, 0, 11, 8, -8, -10, -9, 17, 2, -1, 13, 10, 3, -24, -86, -72, -47, -7, -22, -61, -70, -55, -52, -61, -75, -87, -105, -102, -91, -56, -25, -11, -16, 8, 6, -10, -30, -34, 20, 17, -3, -47, -61, 8, 35, 48, 12, 35, 3, -19, -29, -19, 19, 18, -21, 19, -23, -55, -50, 20, 38, 14, -8, 8, -38, -70, -57, -16, -44, -31, 67, 63, 69, 9, 46, 9, 16, -29, -17, -6, 10, 62, 24, 17, -10, -26, -4, 71, 32, -11, 15, -1, -6, 14, -46, -29, -23, 18, 73, 87, 65, 57, 35, 18, 8, -14, -30, -25, 12, 10, 23, -9, -19, 1, 71, 97, 54, -11, 7, 2, 18, 7, -84, -15, -31, 25, 73, 91, 68, 70, 25, -12, -43, -17, -26, -4, -45, 3, -39, -20, -61, -40, 29, 19, 25, 15, -8, -24, -20, -14, -61, -43, -7, 11, 65, 47, 56, 31, -17, -18, -19, -36, -17, -3, -40, 7, 18, -25, -64, -44, 31, 4, -3, 23, -15, -9, -17, 7, -37, -22, 28, 61, 39, 27, 58, -5, 8, 10, -34, -42, -78, -45, -27, -12, -25, -51, -51, -72, -13, 43, 29, -2, 15, -37, -33, -37, -2, -26, -12, 40, 53, 28, 28, -14, -10, -7, 2, -50, -40, -9, -36, -38, -10, -48, -15, -30, -15, 43, 23, 10, -5, -48, -40, -57, 17, 21, 13, 61, 47, 24, 9, 7, 12, 1, 16, 16, 19, 18, 18, 23, -4, 4, -12, -36, -36, 13, 9, 27, -58, -65, -38, -33, 33, 92, 62, 54, 94, 61, 43, -5, 7, 38, 67, 47, 29, 42, 34, 41, 11, 50, 9, -21, -58, 20, 31, 21, 8, -33, -38, 31, 73, 114, 66, 42, 63, 94, 40, -27, 0, 37, 87, 51, 42, -1, -5, 52, 43, 34, 3, -6, -44, 7, 56, 6, -4, -38, -51, 36, 98, 86, 88, 40, 47, 36, 2, 4, -24, 2, 47, 44, 41, 10, 22, 45, 51, 14, 20, -17, -50, 14, 64, 11, 31, -23, -71, 64, 87, 98, 73, 28, 27, -12, 12, 3, -17, -2, 26, 19, 20, 7, 11, 48, 45, -13, -14, 13, -7, 11, 7, 35, 21, -26, 55, 63, 92, 58, 11, -2, 12, -24, 11, 0, 0, 44, 38, 91, 56, 20, 2, 16, -2, 10, 20, 29, -17, 1, 21, 31, 13, -4, 76, 98, 53, -6, -28, -32, -37, -21, 22, 7, 35, 25, 91, 143, 98, 19, -15, 14, 8, 36, 47, 44, 13, 36, 13, -9, -13, -18, 89, 88, 42, -57, -93, -65, -73, -29, -28, 31, 27, 70, 141, 136, 99, 25, 24, 29, 33, 66, 64, 72, 69, 39, -5, -17, -14, -39, 61, 81, 44, -54, -85, -59, -44, -49, -40, -3, -12, 37, 96, 145, 88, 41, 85, 48, 42, 66, 59, 23, 89, 40, -49, -35, -36, -7, 62, 81, 40, -21, -47, -41, -45, -77, -58, -71, -68, -55, 31, 106, 75, 81, 42, 40, 46, 79, 80, 71, 73, 20, 6, -63, -38, 25, 51, 81, 54, -47, -45, -35, -45, -62, -65, -92, -96, -64, -12, 74, 65, 38, 22, 35, -2, 45, 71, 101, 72, 30, 16, -62, -14, 27, 66, 40, -3, -17, -52, -62, -88, -77, -121, -120, -139, -83, -55, 19, 9, 48, 34, 27, 3, 36, 0, 80, 57, -6, -28, -27, 12, 50, 98, 101, 63, 48, -29, -74, -78, -70, -118, -93, -118, -121, -50, -39, 38, 25, -10, -4, 13, 47, 26, 61, 53, -18, -18, 12, 6, 32, 61, 71, 66, 49, 18, -13, -1, -10, -48, -76, -83, -83, -60, -43, 16, -19, -14, -3, -8, 45, 16, 37, 38, 17, 7, -14, -7, 40, 45, 74, 103, 78, 77, 46, 36, -12, -38, -66, -77, -110, -60, -27, -10, 4, 28, 20, 19, -43, -28, 26, 32, -40, -11, 13, -4, 20, 32, 34, 80, 92, 53, 61, 14, -16, -39, -41, -57, -59, -53, -41, -1, 7, 37, 34, 31, 45, 10, 37, 15, -34, -30, 18, -15, 1, 4, -1, -28, 3, 24, 28, 57, 64, -2, 17, 36, 26, -15, -33, -6, 15, 41, 5, 44, 12, 7, 9, -20, -38, 6, 20, 11, 12, 9, 6, 19, -4, 13, 31, 38, 41, 61, -42, -61, 0, 13, -14, 20, -5, 28, 15, 18, 20, 0, -17, 17, -2, -8, -19, 15, -7, 10, 9, 17, 5, 8, -14, 14, 5, -12, -2, 13, 12, -26, 11, 12, -2, 20, 13, 13, -8, 1, -4, 19, -3, -12, 6, -14, -843, -20, 15, 13, 9, -31, -16, 18, -6, 0, -25, -59, -8, 27, 0, -53, 10, -29, -44, -28, -5, -25, -14, -49, -29, 9, 4, -3, 7, 12, 8, 6, 8, 57, -17, 21, 15, -66, -8, 10, -6, -19, -14, -31, -3, 15, 44, 30, 19, 38, 59, 17, 53, -4, -20, -6, -7, -6, 6, -16, -44, -37, -22, -23, 20, -26, -11, -38, -47, 6, -13, -15, -17, -9, 29, 38, 22, 27, 28, 26, -26, -36, 2, 16, 9, 2, -28, 24, -15, 5, 11, 6, 43, 9, -16, -60, 16, -24, -7, 4, 1, -17, -13, 29, 19, 40, 1, -43, 24, -5, 9, -21, 21, -14, -23, 26, 1, 25, 8, 10, 3, 8, -27, -39, -20, -49, -31, 3, 19, 16, -20, -20, 41, 44, 3, 17, 56, 79, 22, -7, 3, 1, -38, 54, 35, 3, -19, 3, -38, -26, -38, -58, -3, -16, -23, -17, 12, 45, 10, -16, -6, 28, 33, 17, 70, 83, 27, -1, 1, -19, -12, 30, 7, 14, -7, -1, 16, -2, 9, -1, 14, 45, 21, 38, 16, 5, 11, 16, 24, 23, 55, 36, 34, 41, 54, 5, -2, -10, 33, 25, 52, 25, 9, 39, 43, 1, 16, -1, 49, 45, 55, 13, 1, 9, 38, 33, 67, 50, 22, 14, 28, 23, -4, 0, -5, 10, 34, 6, 12, 34, 15, -2, -45, 19, 33, 27, 77, 64, 25, 1, 4, 26, 29, 38, 0, -13, 11, -6, 20, 35, -34, -58, -8, 15, 7, -13, 24, 29, -11, -32, -46, 41, 46, 50, 55, 20, 3, 4, 26, 55, 22, -25, 1, -35, -1, -14, 26, 105, -24, 8, -41, -2, 74, 30, 43, -33, -49, -18, 11, 75, 77, 71, 61, 27, 7, 35, 79, 99, 10, -36, -16, -25, -17, -61, -5, 76, -15, 13, -4, -9, 90, 52, 9, -33, 3, -8, 23, 50, 74, 94, 77, 47, 15, 76, 115, 135, 57, -17, -54, -21, -11, -61, -8, 27, -11, 25, 9, 46, 78, 18, -26, -28, 10, -2, 15, 85, 52, 87, 109, 33, 64, 80, 97, 58, -4, -43, -34, -35, -62, -16, 15, 24, -30, 17, 1, 52, 62, 17, -79, -76, -49, -9, 27, 112, 78, 84, 83, 61, 39, 81, 60, 31, -35, -76, -44, -53, -28, -66, 21, 4, -68, -18, -25, 17, 28, -34, -43, -9, -28, -32, 9, 76, 65, 88, 64, 61, 45, 82, 36, -24, -69, -80, -69, -51, -36, -7, 1, -5, -63, -45, 7, 6, -17, 3, -32, -45, -45, -62, -30, 20, 13, 22, -8, 23, 15, 28, 12, -16, -25, -45, -37, -64, -19, -3, 13, -38, -71, -74, -20, -28, 15, -16, -31, -32, -76, -101, -98, -68, -51, -61, -32, -64, -43, -23, 8, 5, -4, -37, -20, -1, -11, 12, -14, -52, -124, -74, -28, 28, 17, -38, -52, -14, -36, -67, -76, -82, -69, -35, -74, -60, -38, -43, -9, 5, -21, -49, -21, -43, -38, -63, -34, -56, -76, -29, -48, -27, 49, -16, -41, 1, -16, -27, -51, -35, -45, -52, -47, -21, -20, -15, -16, -7, 1, -31, -33, -55, -62, -51, -54, -39, -43, -50, -17, 7, 64, 23, 15, -7, 11, -19, -14, 1, -15, 14, 39, 23, 40, 53, 24, 35, 7, -46, -36, -25, -22, -48, -13, -57, -30, -49, -12, -27, 30, 68, 46, 34, 8, 51, 45, 27, 45, 52, 77, 93, 54, 44, 23, 42, 3, -20, 12, -46, -32, -64, -24, -26, -15, -29, 14, 2, 29, 49, 41, 26, 16, 46, 63, 64, 66, 70, 83, 69, 15, 33, 29, 47, 50, 66, 10, -27, -24, -92, -53, -3, -5, -3, 16, 9, 20, 55, 18, 47, 58, 41, 89, 44, 64, 39, 48, 37, 16, 37, 68, 43, 21, -17, -8, -1, -18, -6, -5, 29, -19, -2, -2, 30, 24, 43, 13, 4, 32, 18, -9, -3, -25, -10, 10, 12, 58, 53, 39, 3, -19, -24, -2, -29, -45, -28, -25, -44, -2, -9, -14, -16, -20, -4, 4, 2, 4, -11, -7, -29, 12, 0, -12, -4, -8, -21, -11, -24, -36, -57, -69, -54, -27, 5, -39, -19, -22, -17, 4, 5, -15, 14, -7, -22, -60, -49, -19, -39, 11, -11, -36, 3, -7, 19, 3, 1, -41, 17, -26, -35, -36, -25, -37, -13, -17, 15, -17, 6, -4, -2, -17, -6, -37, -28, -59, -35, -28, -32, -9, -50, 6, -45, -56, -82, -31, -52, -33, -19, -4, -12, 13, 13, -15, 1, -20, -12, 5, 17, -14, 16, -3, 4, 13, 8, -6, -15, -3, 6, -1, 11, 1, 1, 10, -8, 17, -3, 13, 14, -4, -2, 1, 1, 14, 817, -19, -9, -6, -7, 30, -16, -35, -12, -48, -64, -56, -52, -95, -151, -36, -41, -56, -17, -62, -33, -49, -12, 27, -4, -21, -15, -3, -19, -14, 13, -13, -36, -34, -8, -28, -61, -83, -87, -97, -52, -103, -162, -99, -78, -91, -119, -143, -150, -140, -122, -76, -57, 13, 14, 14, -2, 6, 24, -20, -6, -19, -7, 11, -59, -55, -62, -35, 9, -28, -77, -56, -66, -59, -60, -120, -135, -146, -87, -84, -80, -9, 1, -10, -15, -6, -12, 7, 4, -31, -12, -15, -81, -52, -77, -59, -21, -17, 8, -8, -24, -50, -75, -39, -123, -116, -79, -70, -55, 17, -25, -8, -7, 7, 19, 7, -56, -64, -56, -31, -77, -88, -88, -49, 3, 9, -12, -7, -4, -15, 15, -13, -47, -55, -85, -103, -63, -55, -19, -16, -11, 14, 56, -2, -60, -79, -43, -44, -52, -31, -62, -17, -6, 15, -18, 36, 34, 53, 14, 26, -44, -42, -82, -76, -58, -21, -37, -5, 0, 15, 57, -29, -82, -59, -14, -26, -53, -39, -58, -13, 4, 3, 12, 26, 57, 84, 44, 10, -22, -34, -54, -48, -39, 43, -50, 9, 2, -18, -23, -68, -85, -96, -61, -67, -52, -37, -29, -26, -31, 19, 15, 58, 88, 85, 55, 28, -7, -16, -35, 8, -30, 17, 36, 20, 19, -10, -43, -99, -47, -26, -43, -48, -17, -38, -3, 7, -15, 23, 39, 68, 60, 65, 48, 5, -19, -31, 22, 3, 24, 18, 47, 54, -18, -32, -63, -53, -11, -27, -66, 5, -28, 10, 45, -13, 26, 25, 18, 30, 48, 3, -20, -6, -5, -7, 4, 39, 53, -13, -12, -2, -19, 8, -52, 6, 22, 8, -9, -5, 25, 26, 59, 41, 15, 2, -12, -4, 1, -3, -12, -4, -7, -20, 10, 45, 57, -2, 18, 3, -7, -5, -21, 55, 42, 26, -8, 30, 25, 58, 60, 45, -10, 6, -17, -17, 8, 3, 20, 20, 18, 24, -15, 18, 6, 84, 7, 4, -30, -29, -23, 30, 46, 36, 29, 40, 13, 20, 29, 33, 6, -22, -52, -33, 5, 21, 43, 57, 35, 61, 39, -3, -26, 26, 25, -8, 7, -57, -86, 23, 79, 69, 30, 5, 17, 37, 1, 39, -17, -46, -51, -46, 53, 82, 106, 88, 50, 9, -7, 25, -39, 25, 38, 27, 9, -39, -23, 33, 65, 46, 6, 15, 6, 16, 3, 17, -21, -38, -77, -24, 75, 81, 76, 45, -2, -34, -7, -26, -76, 18, 23, 43, 10, -59, -29, 6, 33, -5, 23, 17, -11, 3, 6, 3, -24, -26, -54, 40, 84, 83, 64, -4, -21, -67, -59, -77, -93, 29, 3, 14, 13, -62, -47, -42, 1, -10, 15, -3, -18, 20, 2, 13, 29, -14, -53, -17, 23, 39, 9, -5, -79, -63, -102, -49, -52, 2, 20, 43, 9, -48, 4, 7, 52, 12, 22, 1, 9, 36, 39, 54, 30, -16, -70, 17, 25, 16, -3, -4, -45, -66, -99, -35, -23, 17, 37, 21, 13, -17, -47, 60, 55, 25, -25, 32, 12, 16, -7, -9, -10, -103, -70, -46, 1, -4, -15, 6, -18, -65, -118, -76, 2, -63, 2, 16, 10, -14, -46, 64, 15, 24, -13, -28, -13, -62, -61, -57, -85, -98, -111, -54, -13, -1, 8, 31, -8, -28, -93, -24, 5, -26, 9, -5, 19, 34, 5, 28, 19, 23, -10, -52, -103, -104, -108, -108, -122, -136, -85, -65, -24, 12, -2, 28, 4, -4, -62, 25, 1, -46, 7, 13, -15, 10, 25, -13, 71, 76, 32, -47, -90, -75, -106, -98, -112, -104, -89, -63, -26, -40, -18, 7, -10, -58, -69, 11, -2, -49, 22, 14, -1, 28, 31, -19, 62, 119, 95, 38, -4, 16, -11, 3, 11, -41, -17, -39, -43, -21, 6, 5, -30, -28, -60, -1, 4, -23, -38, 13, -6, 28, -22, -7, 42, 68, 65, 91, 101, 102, 58, 55, 32, 24, 30, -17, -27, -9, -5, -22, -58, -6, -30, -4, 13, -21, -52, -15, 12, -12, 28, -24, 13, -20, 25, 53, 60, 68, 69, 65, 58, 42, 47, 10, 17, 38, 12, 36, 55, 36, 30, 16, 26, -7, -17, 0, -12, -5, 14, -34, -10, 37, 54, 51, 26, 76, 38, 33, -32, -2, -5, -8, 25, 7, 28, 30, 72, 58, 64, 23, 15, 13, -19, -9, 6, 19, -18, 11, 10, 19, 43, 48, 52, 19, 46, 6, 1, -44, -56, 32, 45, 11, 40, 45, 31, 39, 45, 4, 22, -4, -15, -21, 19, 2, 6, 16, -20, 18, -7, 1, 0, -19, -7, 1, -12, -14, -30, 16, 13, 1, -16, 20, -4, -17, 20, 17, -19, 0, -19, -19, -10, 456, 12, -14, -5, -20, -37, -9, -15, 7, -14, -28, -41, -24, 31, 14, -38, 8, -6, -31, -15, -19, -1, -1, -32, -19, 2, 0, 9, 15, -4, 6, -27, 11, 13, -28, -12, -17, -46, -1, 2, -29, -73, 24, 2, 26, 0, 27, 37, 24, 19, 59, 10, 70, 19, 5, 17, 1, 9, -41, -5, -52, -12, -34, -8, -2, -22, -30, -47, -45, -25, 11, 7, -23, -22, 4, -9, 20, 0, 25, -35, -61, -44, 37, 19, 1, -11, -46, -67, -55, 45, 23, 12, 19, 9, -35, -38, -29, -44, -20, 12, -4, 21, 29, 2, -7, 11, -26, -46, -50, -12, 3, -5, -15, -17, -42, -29, -64, -8, 36, 19, -25, 12, 4, -34, -11, -24, -6, -18, -13, -38, -38, -42, 0, -13, -25, -16, 0, 42, 85, -8, 1, 16, -47, -42, -74, -61, -16, -23, -35, -33, -11, -7, -6, -24, -7, -13, -46, -46, -29, -68, -38, -12, -1, -6, 5, 42, 26, 16, 16, -22, -71, -55, -95, -96, -44, -42, -37, -46, -60, -19, 0, -32, -45, -35, -67, -44, -60, -29, -40, -29, -3, 6, 23, 40, 11, 31, -20, -25, -43, 2, -53, -71, -69, -25, -25, -41, -49, -34, -34, -74, -70, -73, -116, -103, -67, -77, -85, -58, -15, 7, 5, 74, -1, 21, 15, 2, -49, -29, -88, -44, -28, -39, -38, -26, -42, -52, -52, -94, -71, -24, -31, -41, -2, -32, -34, -57, -7, -1, -10, 78, -24, -40, 11, -16, -41, -51, -57, -45, -43, -65, -23, -26, -52, -32, -45, -31, 6, 77, 53, 51, 10, 33, -20, -19, 14, -6, -9, 41, 13, -7, 2, -59, -42, -70, -30, -27, -56, -58, -25, -39, -14, -29, -4, 15, 49, 113, 88, 46, 12, 8, -12, 8, 26, 26, 38, 35, 8, 19, -1, -36, -62, -34, -48, -12, -46, -57, -32, -13, 30, 5, 31, 28, 70, 115, 81, 61, 44, 31, 12, 30, 53, 39, 52, 43, 1, 19, -3, -19, -35, 0, -98, -9, 26, -8, 14, 74, 73, 47, 44, 43, 100, 132, 107, 112, 66, 42, 70, 17, 39, 47, 47, 27, -49, 35, 2, -49, -30, 15, -64, -37, 30, 54, 84, 99, 65, 68, 70, 59, 94, 152, 98, 87, 20, 0, 24, 6, 25, 19, 52, 44, -108, -9, -38, -3, -57, -18, -49, 23, 35, 81, 105, 90, 49, 31, 65, 118, 126, 101, 49, 6, -30, -37, -10, -26, -17, -1, 86, 25, -89, -18, -17, -48, -42, -62, 3, 55, 44, 59, 54, 61, -4, 3, 66, 103, 93, 25, -63, -65, -93, -41, -50, -54, 5, 20, 19, -18, -70, -65, -12, -10, -18, 16, 46, 31, 26, 40, 27, 6, -13, 5, 50, 70, 18, -85, -100, -85, -64, -41, -51, -36, 0, -8, -25, -17, -81, -51, -31, 9, -53, -54, -17, -11, -20, -4, -7, -9, -4, 24, 40, 3, -96, -112, -92, -50, -50, -26, -40, -38, -21, -18, -20, -57, -89, -17, -5, -45, 56, -25, -38, -21, 1, 25, -17, 9, 5, -16, -21, -54, -74, -64, -60, -6, -38, -53, -43, -30, -22, -35, -84, -19, -47, -52, -17, 31, 59, 13, 15, -28, 9, 17, -20, 41, 25, -3, 11, -19, -32, -15, -19, -15, -25, -6, -49, -25, -9, -9, -7, 12, -32, -77, -18, -17, 4, 17, -3, -3, -17, -15, -7, 10, 14, -11, -6, 23, -19, 6, 1, -23, 22, -27, -23, -25, -13, -4, -12, -17, -29, -56, 18, 23, 4, 34, -4, 19, -37, -20, 12, 21, 6, 1, 5, 22, 14, 21, 19, 7, 29, 25, 44, 62, -1, -14, -21, 10, -9, -8, 6, 3, 36, 16, 19, -25, 1, -1, -13, -34, -40, -32, -4, 29, -9, 9, 52, 58, -11, -11, 15, 66, 62, 22, 22, 18, 3, 14, -4, 27, 49, 1, 9, -44, -28, -1, 21, -25, -26, -24, 33, 17, 25, 10, 16, -9, 18, 24, 36, -10, 1, 1, 16, 17, -9, -14, 8, -15, -32, -17, -2, 18, 12, -18, -13, -56, -61, -26, -72, -33, -68, -44, -92, -72, -68, -127, -92, -64, -69, -18, -47, -22, -25, -20, -1, -12, 4, -55, -37, -41, -34, -34, -37, -91, -51, -59, -98, -87, -56, -71, -53, -58, -93, -72, -83, -72, -33, -20, -56, -17, -22, -5, 18, -8, 17, 4, 12, -14, -42, -18, -17, -42, -31, -50, -60, -6, 23, -3, -47, -33, -41, -36, -49, -31, -53, -16, 12, 16, -11, -20, 15, -5, 11, -14, -16, 15, 4, 16, 9, 4, 0, -5, -9, 11, 10, 0, -14, 1, -20, 3, 0, 2, -10, -11, 12, -9, 16, -17, -9, -1228, 9, 3, 18, 6, 4, 37, 35, 61, 32, 63, 107, 78, 83, 118, 38, 28, 9, 32, 56, 31, 42, 38, -3, 7, 5, -2, 15, -11, 10, -18, 3, -6, 39, 47, 43, 66, 70, 73, 53, 46, 102, 142, 82, 37, 62, 111, 111, 117, 118, 125, 89, 37, 16, -17, 18, -1, 16, -13, 23, -25, -46, -27, 31, 56, 32, 16, 9, 39, 33, 73, 13, -3, 31, 16, -26, 5, 17, 15, 38, 60, -31, -7, -12, 13, -17, -28, -9, 19, 14, -11, 10, 6, 12, 3, -1, 32, 14, -12, 7, -39, -15, -30, -59, -50, -35, -49, 6, 6, -87, 1, -2, 4, -9, -96, -44, 14, 12, 23, -19, -17, -1, 17, 12, 6, 5, 10, 24, 14, 4, -58, -52, -38, -98, -92, -78, -71, -68, -41, -1, 18, -9, -47, -76, -23, -44, -46, -28, -38, -67, -21, -47, 0, -4, 18, 23, 10, 10, -16, -43, -13, -93, -83, -113, -98, -65, -27, -21, -5, 1, -10, -13, -2, -22, -70, -49, -58, -16, -29, -31, 15, -9, -31, -9, -15, -2, -16, -22, -22, -65, -82, -96, -110, -89, -29, -14, -12, -3, -15, 18, 15, -24, -36, -62, -28, 2, -39, -41, -23, -48, -32, -30, -5, -9, 37, 9, 1, -61, -146, -160, -176, -104, -23, 5, 7, -31, 21, -47, -58, -16, -43, -50, -20, -5, -11, 2, -29, -29, -34, -61, -35, 7, 74, 39, -23, -50, -123, -130, -112, -67, 17, 19, 14, -14, 17, -4, -54, -34, -33, -24, -5, -5, -16, -15, -17, -21, -52, -51, -17, 40, 73, 22, -46, -80, -106, -91, -112, -75, 9, -21, 41, 54, 44, 23, 4, -37, -27, -48, -21, -42, -18, 18, -10, -22, -15, -12, 37, 29, 31, -14, -60, -113, -84, -69, -40, -51, 0, -19, 16, 75, 39, -23, -10, 19, -4, -10, -5, -13, 17, 18, 30, -26, -57, -11, 1, 9, -23, -58, -71, -77, -80, -44, -6, -67, -41, -2, 6, 48, 32, 12, 30, 32, 29, -27, 30, 8, 12, 21, 4, -7, -38, -19, -26, -28, -43, -95, -104, -96, -78, -56, -20, -27, -31, -34, -21, 51, 97, 27, -23, 18, 12, 33, -16, -5, 28, 10, 2, -24, -29, -49, -69, -33, -51, -108, -82, -58, -64, -46, 36, 7, 31, 31, -27, 40, 64, 40, -14, 7, 57, 7, 5, -15, 6, 39, 39, 8, -32, -58, -84, -52, -53, -68, -49, -14, 14, 15, 75, 48, 47, 46, -5, 40, -2, -3, -11, 6, 14, -1, 3, 19, 47, 45, 26, 14, -37, -70, -100, -73, -65, -24, -2, 19, 72, 79, 61, 40, 43, 19, -20, 18, 26, -33, -24, -26, 13, -4, 26, -12, 39, 25, -3, -6, 5, 3, 10, 7, 21, 31, 39, 96, 98, 73, 25, 43, 45, 43, 19, 49, -4, -41, -57, -43, -18, -26, -2, 9, 23, 10, -11, -46, 31, 23, 21, 34, 19, 58, 44, 74, 91, 77, 19, 54, 45, 8, 11, 26, 43, -18, -59, -73, -43, -38, -24, 22, 20, 1, -33, 3, 16, 27, 32, 27, 58, 55, 45, 33, 38, 22, 9, 20, 6, 49, -2, 19, 28, -39, -95, -59, -62, -30, -38, -12, 3, 4, 11, 15, 40, 18, 14, 26, 44, 23, 59, 22, 20, 0, 20, 5, 11, 27, -23, -9, 5, -39, -107, -107, -78, -51, -75, -40, -24, -20, 11, 45, 51, 26, 23, 8, 6, 22, 27, 0, 13, -72, -1, 47, 41, -14, -19, 6, 25, 24, -77, -91, -86, -45, -66, -57, -10, 28, 25, 61, 48, 61, 25, 32, 36, 28, -11, -40, -32, -54, -24, 68, -16, 5, -6, -20, 44, 45, -7, -54, -91, -57, -82, -84, -57, -17, -20, -24, 25, 61, 64, 67, -36, -28, 1, -63, -49, -22, -43, -5, -21, 17, 10, 21, 56, 24, -1, -12, -35, -26, 0, -28, -70, -77, -72, -75, -76, -62, -31, -43, -101, -92, -32, -41, -60, -38, -45, 10, -15, -12, -19, 13, -4, 21, 7, 47, -8, -15, -84, -66, -38, -83, -118, -162, -147, -138, -135, -117, -152, -101, -104, -106, -68, -31, -4, 15, 3, 20, -7, -11, 14, 3, 40, -45, -43, -42, -87, -89, -14, -92, -90, -155, -163, -97, -69, -44, -56, -37, -76, -53, -14, -2, -7, -7, -8, 3, -5, 10, -13, -20, -19, -9, -38, -63, -33, -33, -66, 0, 26, -13, -38, -46, -25, -41, -32, -17, -24, -46, -41, 12, 15, 9, 20, 21, -18, -2, -7, -7, -1, -6, -12, 15, -1, 10, 9, 16, -20, -14, -2, 7, 9, 15, 20, 20, -6, 11, -5, -7, -5, -15, -21, 12, -2, -298, 5, -18, 6, -1, 49, 56, 21, 28, 14, 22, 47, 11, -37, -5, 38, -13, -15, 47, 13, 35, 20, 25, 40, -4, 7, -13, 2, -11, 10, 15, 5, 1, -31, 29, -31, -17, 44, 31, 45, 19, -26, -40, 3, -26, 15, 23, -20, -26, -65, -46, -67, -69, 2, 12, -18, -12, 2, 34, 1, 49, -19, -8, -27, -29, 37, 60, 56, 45, 38, -8, 31, 26, 31, 7, 9, -19, -29, -7, 15, 0, -19, -41, -12, -11, -3, 30, 22, 37, -47, -47, 2, -21, -1, 24, 41, 46, 55, 49, 54, 64, 27, 27, 3, -20, -40, -12, -16, 15, 50, 31, -11, -13, 19, -49, 39, 47, -27, -7, -28, -16, -3, -16, 8, 33, 53, 31, 70, 47, 78, 61, 53, -4, 18, -24, -28, 26, 51, 37, 4, 0, 12, -35, 60, 37, 48, 25, 22, 29, 10, -2, 15, 32, -14, 21, -10, 15, 24, 34, 9, 41, 20, 34, 11, 45, 30, 20, -18, 7, 19, 44, 66, 43, 56, 32, 37, 40, 31, 21, 3, -35, -16, -33, -40, -31, 11, -27, -20, 26, 38, 64, 25, 84, 39, 41, -5, -15, 11, 1, 12, 54, 46, 46, 36, 40, 17, 6, -20, -42, -20, -27, 16, -17, -19, -29, 2, 47, 32, 72, 100, 96, 112, 21, 14, 20, 8, 30, 22, 45, 52, 32, 47, 30, 56, 39, 15, -27, 1, -18, 40, 1, -52, -26, -41, 25, 18, 87, 93, 150, 68, 34, 51, -7, 2, -20, 0, 60, 25, 59, 25, 46, 43, 1, 1, 28, -7, -4, -42, -50, -16, -29, -16, -6, -12, 77, 123, 112, 83, 6, -1, 30, 65, 31, 22, 23, 46, 29, 24, 53, 16, 19, 35, 17, -51, -59, -86, -54, -44, -58, -60, -55, -67, 11, 128, 144, 104, -12, 10, 2, 34, 57, 33, 39, 15, 4, 2, 39, 25, -18, 7, -33, -88, -94, -59, -48, -67, -50, -53, -112, -87, -9, 85, 128, 100, 15, 5, 17, 16, 7, 27, 59, -11, -41, -27, -8, 6, -13, -75, -70, -71, -68, -58, -21, -39, -37, -43, -80, -93, -26, 28, 58, 67, -21, -16, 7, 23, 39, -7, 24, -21, -72, -79, -12, -1, -49, -25, -74, -44, -43, -50, -36, -32, -47, -68, -61, -64, -56, -30, -27, 56, 57, -17, 25, -1, 38, -31, -10, -70, -41, -55, -22, 3, -13, -33, -51, -55, -29, -21, -10, -39, -41, -53, -58, -55, -91, -45, -105, 45, 50, -3, -4, -23, 63, 37, -13, -74, -70, -60, 8, -4, -45, -16, -40, -44, 3, 6, 12, 2, -51, -28, -28, -24, -75, -58, -61, 65, 32, 29, -13, -34, 68, 83, 37, -30, -20, -24, -8, -5, 2, 3, 10, 40, 58, 30, 29, 42, 1, -33, -10, 2, 1, 10, 25, 93, 86, 70, 35, 31, 87, 83, 56, 25, 30, 18, 33, 24, 53, 53, 81, 51, 71, 29, 28, 39, 37, 49, 41, 41, 50, 49, 29, 71, 83, 43, 20, 44, 93, 96, 88, 89, 41, 51, 39, 13, 69, 81, 72, 55, 36, 17, 52, 47, 62, 48, 55, 41, 42, 55, 7, 54, 53, 25, 20, 25, 51, 22, 43, 78, 63, 38, 33, 15, 37, 72, 72, 51, 43, 26, 41, 27, 69, 39, 39, 75, 48, 42, 3, 55, 31, 63, 25, -22, -7, -10, -4, 23, 21, 2, -27, -6, 3, 20, 29, 22, 39, 19, 51, 40, 38, 51, 60, 51, 79, 23, -14, 51, 61, 37, -3, -14, 23, -15, -33, 17, 23, 14, -12, -1, -12, 5, 24, 21, 14, 36, 40, 41, 53, -1, 21, 12, 18, -35, -13, 70, 41, 33, 1, -28, 10, 1, -50, -31, 30, -2, -3, -18, -15, -3, 52, 57, 33, 32, 14, 72, 7, 19, 1, 12, -15, -53, -24, 46, 3, 9, 20, 0, 34, 38, 10, -63, -39, -36, -22, -41, -32, -23, -4, 40, 44, 23, 34, 63, 9, 32, -15, 4, -32, -42, -15, 45, 4, -10, -20, 3, 16, 16, -25, -48, -66, -24, 27, -29, -1, 10, 8, -25, 8, -11, 17, -17, -9, -5, -28, -13, -40, -21, 1, 8, 18, -12, 7, -3, 4, 7, 17, -16, -14, -35, -15, -23, 0, -14, -32, -72, -73, -73, -49, -66, -50, -34, -2, -17, -20, 0, 2, 26, 9, -15, 10, 16, 4, -17, 18, 0, -28, -37, -16, -48, -25, 10, 5, -36, -32, 11, 16, 13, -21, -23, -13, -10, -1, 17, -13, -20, -9, 0, 17, -9, 13, -3, -3, 4, 17, 1, -2, 6, -6, -16, 13, 11, 22, 11, 6, -9, -2, 20, -11, -18, 18, -11, -9, 3, 6, 19, 4, 1272, -8, -14, -16, 3, -16, 16, 1, -17, 18, -20, -49, -14, -4, -6, -54, -56, -25, -19, -39, -22, -31, -42, -16, -13, -8, 17, 5, 5, -3, 4, -7, 5, 27, -14, 14, -11, -69, -7, 1, -81, -77, -17, -25, -6, 13, 1, -12, -21, 22, 31, 41, 47, 18, -14, -20, -12, 2, -29, -18, -6, 2, 30, 66, 50, 12, 9, 9, 14, 26, 14, 14, -7, -37, -16, -35, -45, -54, -31, -31, -78, -25, 3, 0, 16, 16, -43, -74, -63, 24, 24, 42, 77, 54, -7, -52, 31, -21, -35, -31, -8, 2, 2, -37, -1, -72, -56, -100, -130, -51, -12, 15, -6, -17, -29, -21, -46, -48, 1, 14, 4, 12, 4, -21, -14, -25, -20, -29, -37, -75, -61, -44, -37, -55, -44, -24, -41, 19, -28, -13, -2, 3, 8, 8, -48, -65, -64, -24, -5, -15, -21, -28, -42, -57, -24, -25, -59, -65, -64, -96, -39, -19, -17, -29, -3, -8, -70, -21, 19, -2, -44, -33, -47, -77, -14, 5, -13, -19, -37, -7, -64, -55, -74, -86, -86, -69, -47, -29, -45, -27, 5, 8, -43, -87, -41, -21, -10, 11, -33, -55, -32, -33, 15, -2, -16, -42, -24, -35, -41, -72, -67, -45, -47, -20, 8, -2, -41, -16, 3, 7, -36, -69, -29, 5, 16, -24, -43, -79, -31, 27, 32, -27, -20, -28, -15, -43, -23, -45, -20, 14, 25, 36, 60, 72, 24, -18, 28, 59, 26, -62, -48, -16, 6, -35, -1, -26, 2, 1, -22, 3, 13, -21, -10, -3, 5, 36, 71, 66, 91, 60, 60, 65, 43, 22, 97, 57, 26, -17, -7, -7, -24, -42, -20, -28, 15, 38, 21, 23, 13, 8, 20, 21, 40, 65, 94, 87, 74, 60, 57, 85, 93, 67, 97, 45, 23, -22, -16, -20, -7, -48, -80, 3, -21, 60, 34, -15, -21, -6, 26, 46, 54, 74, 66, 28, 31, 59, 56, 73, 80, 62, 56, 20, 25, -30, -71, -3, -6, -25, -77, 33, 19, 62, 61, 3, 8, 32, 13, 28, 57, 45, 72, 81, 73, 57, 71, 67, 56, 25, 21, 9, 19, 0, -17, -31, -10, -34, -42, 24, 29, 52, 56, 25, 11, 37, -6, 21, 37, 56, 27, 62, 48, 62, 13, 41, 14, 20, 16, 30, 44, 26, -22, 3, 10, 22, 8, -14, 38, 57, 94, 41, 13, 7, -11, 15, 58, 78, 70, 49, 9, 26, -22, 14, 27, 34, 21, 44, 69, 53, 2, 25, 19, -6, 36, 13, 19, 48, 77, 71, 13, 26, 1, 30, 99, 99, 140, 81, 42, 2, 5, 33, 34, 70, 46, 85, 81, 81, 19, -6, -14, 35, -31, -7, 13, 31, 38, 29, 9, 1, 17, 46, 79, 124, 134, 91, 58, 20, 51, 56, 72, 61, 72, 41, 52, 19, -18, -33, -20, -26, -8, -27, 25, 57, 5, 11, -1, 16, -10, -25, -4, 55, 53, 47, 60, 60, 50, 65, 55, 78, 29, 26, 54, -18, -51, -23, -18, -8, 48, -2, 17, 21, -13, 13, -16, -5, -22, -39, -49, -78, -67, -19, -2, 38, 56, 23, 16, 3, 56, 80, 24, -25, -26, -40, -35, 10, 24, 38, 12, -8, 15, 12, 7, -29, -63, -37, -62, -104, -83, -47, -31, -7, -13, 5, -27, -9, 23, 24, -27, -25, -42, -65, -41, -12, -18, -20, 2, -11, 19, -11, -16, -57, -57, -74, -45, -37, -84, -76, -63, -26, -11, -45, -38, -14, -41, -6, -37, -60, -40, -66, -14, 2, -23, 3, -15, 18, -49, -7, -21, -15, -40, -13, -43, -18, -40, -48, -40, -27, -39, -19, -10, -19, -59, -55, -68, -112, -41, 0, -1, 60, 1, -8, 24, -27, -36, -4, 2, -13, -27, -16, -55, -32, -68, -62, -16, -23, -11, -27, -64, -30, -78, -101, -66, -66, 18, -11, 9, 27, -54, -10, 53, 18, -18, 30, 15, 15, -14, 20, 15, -2, 1, -30, -19, -70, -21, -60, -31, -18, -35, -34, -10, -29, -19, 17, 13, 20, -14, 16, 37, 101, 116, 76, 3, 3, 21, -19, -12, 3, -36, -64, -91, -80, -67, -19, -52, -26, -3, -8, 10, -4, -33, 20, -13, 2, -8, 2, -15, -13, 22, 36, 36, 31, 48, 78, 80, 65, 47, -1, 1, 2, -13, -23, -8, 21, -5, 13, 20, -16, 4, 10, -9, -5, 6, -19, 16, -21, 5, 26, 8, 29, 1, 4, -16, 42, 19, 30, 18, -9, 4, -8, 3, 6, -6, 20, 20, -14, 14, -7, -2, 7, 3, -14, 16, 9, 13, -5, 4, -13, 14, -13, 2, 4, -24, 19, 7, 12, -17, -17, -2, 12, -8, -13, -4, -3, 7, 7, -7, 664, 0, -19, -15, -18, -4, -2, -5, -27, -2, 11, -11, 30, 52, 101, 23, 44, 16, 29, 21, 11, 24, 32, -11, 1, 7, 5, 10, -2, -16, 9, 18, -4, 12, 12, 11, 1, -13, 42, 69, 52, 55, 74, 33, 28, 56, 38, 41, 39, 78, 70, 61, 74, 8, -1, 20, -17, 0, -36, -19, -37, -48, -28, -68, -14, -73, -59, -22, -22, 17, 13, -38, 2, 34, 18, 28, -9, 41, 36, 1, -30, 13, 24, 17, 7, 11, -2, -33, -56, -63, -80, -66, -109, -103, -86, -83, -17, 12, 5, 7, 42, 25, 32, -6, 8, 18, 11, 4, -100, -85, -43, 17, -2, -2, -38, -2, -39, -62, -127, -142, -117, -152, -119, -88, -9, 1, 0, 32, 32, -6, 3, 4, 13, 13, 7, 3, -8, -30, -38, 7, -13, -21, -17, 10, -62, -113, -117, -154, -165, -118, -126, -61, -55, -18, 1, 15, 25, 35, 9, -15, -7, 22, 26, -32, -20, -29, -41, -19, -11, -19, -16, -29, -82, -114, -141, -134, -110, -114, -99, -22, -35, -35, -40, -14, -6, 19, 22, -6, -35, 4, -19, -59, -103, -119, -55, 3, 14, -6, 18, -40, -78, -114, -115, -143, -134, -86, -68, 15, 9, -23, -31, 5, -2, -4, 8, -24, -22, -4, -55, -78, -137, -178, -53, -12, 2, -6, 16, -17, -90, -155, -146, -133, -118, -93, -20, 31, 18, -24, -14, 19, 25, -19, -3, -30, -11, -24, -39, -93, -120, -159, -44, -35, -7, 2, -16, -61, -132, -130, -141, -121, -103, -87, -54, 14, -34, 4, 17, 51, 35, 4, 1, 4, -28, -11, -15, -74, -73, -108, -40, -1, -1, -61, -25, -100, -129, -139, -131, -150, -164, -186, -71, -39, -26, 11, 31, 41, 0, 22, 5, 39, 2, 7, 9, -15, -21, -39, -20, -12, 19, -35, -40, -98, -114, -140, -113, -120, -187, -182, -111, -55, 11, 17, 65, 34, -4, -12, 18, 1, -59, -58, -15, 12, -34, 32, -36, 2, -7, -28, -71, -73, -67, -123, -82, -87, -123, -113, -62, -20, 20, 47, 78, 16, -24, -36, -32, 7, -7, -32, -21, -33, -43, 8, 20, 10, 27, -38, -66, -47, -38, -100, -88, -65, -66, -47, -118, -26, 8, 45, 66, 4, -37, -63, -27, -37, -14, -63, -89, -72, -33, -23, -18, 1, 11, -9, -49, 1, -6, -16, -13, -10, 28, -47, -79, -33, 21, 57, 22, -29, -13, -43, -27, 11, -10, -42, -88, -93, -12, -15, -60, -28, -9, -24, 29, 11, 73, 60, 26, 17, 1, -44, -68, 2, 13, 38, 4, -24, -35, 16, 2, 30, -12, -68, -46, -24, 7, -6, -34, -31, 13, 32, 104, 67, 126, 94, 88, 73, -8, -38, -12, -20, 17, 25, 31, 27, 24, 16, 24, 12, -19, -93, -94, -79, -32, -49, -21, -55, 2, 52, 51, 118, 115, 71, 60, 85, 44, 20, 12, -48, -6, 28, 47, 62, 48, 16, 25, -54, -74, -138, -159, -79, -29, -100, -71, 11, -18, -19, 78, 150, 99, 14, 24, 81, 42, 14, 21, -18, -49, -18, 40, 74, 88, 36, -22, -72, -96, -51, -33, -57, -30, -66, -57, -51, -23, 31, 95, 94, 99, 36, 26, 20, 41, 60, 15, -21, -29, -21, 15, 51, 85, 27, -40, -44, -78, -56, 8, -14, -31, 14, -7, -76, -27, 27, 46, 26, 26, 45, 3, -3, 17, 41, 15, -17, -40, -43, -30, -8, 24, 10, -40, -92, -118, -62, -70, -46, -24, -9, 11, -61, -3, 23, 66, 83, 45, 35, 13, -5, 32, 35, -3, -37, -60, -48, -26, -34, 2, -27, -75, -119, -96, -84, -98, -36, -37, -13, 5, -22, 4, -40, 39, 60, 12, -10, -34, -48, -12, -47, -67, -41, -39, -22, 17, 11, -36, -43, -78, -73, -68, -38, -52, -61, -74, 1, 41, 9, 13, -40, 45, 40, 19, 44, -10, -41, -60, -66, -57, -37, -43, -17, -9, -46, -67, -72, -90, -75, -69, -74, -60, -46, -29, 40, 27, -4, -19, -16, -4, 37, -46, -38, 21, -35, -34, -23, 24, -53, -51, -26, -27, -9, -27, -100, -94, -53, -72, -52, -17, -48, -21, -26, 12, -13, -18, -13, -5, -45, -35, -53, -47, -67, -20, -10, -37, -40, -29, 2, -26, 17, -73, -76, -60, -62, -22, -16, 0, 12, -24, -27, 13, 6, 0, -16, -19, 21, -4, -10, -29, -26, -30, -12, -14, -35, -73, -2, 44, -11, -14, -35, -19, 0, -29, 4, 12, -19, 12, 15, -13, 6, 5, 12, 0, -14, 2, -18, 19, 3, 14, -3, 14, 3, -14, -20, 10, 14, -10, -3, -11, 0, -13, 4, 14, -20, 20, 1, -16, 18, -1, -972, 12, 13, -5, -8, -15, -6, 18, 6, 46, 52, 54, 70, 83, 110, 31, 25, 1, -1, 38, 31, 58, 12, 24, -11, 12, 0, -7, 15, 1, 17, 0, 29, 5, 30, 51, 24, 33, 67, 64, 19, 4, 75, 11, 1, 17, 41, 47, 82, 83, 39, 26, 0, -10, 15, -12, 11, 0, 9, 35, -25, -59, -83, -15, 63, 50, 39, 9, -56, -38, 3, -18, -43, -7, 41, 22, 24, 23, 21, 22, -28, -31, 29, 7, 4, 15, 25, 49, 25, -12, -13, 13, 31, 30, 14, -40, -6, -31, -64, -57, -19, -5, 47, 24, 35, -1, -39, -49, -8, -44, 5, 18, -1, 12, -20, -29, -15, -1, 25, 5, -5, 1, 15, -16, -8, -53, -46, -39, -28, -19, 15, 26, 36, 49, 8, -10, -14, -25, 7, -15, 4, -6, -55, -34, -13, -14, 17, -19, -40, -16, -30, -19, -36, -50, -44, -25, 5, 32, 47, 57, 50, 46, 63, 23, -7, 16, 44, 10, 20, -9, 2, -6, -25, -22, -13, -30, -68, -34, 11, -4, 14, -2, 5, 15, -7, 18, 30, 16, 47, 28, 51, 20, -33, 20, 57, -9, -15, -8, 47, 13, 3, 31, 8, -5, -27, -48, -25, -18, 22, -5, 2, 23, 3, 11, 35, -25, 24, 31, 6, 36, -35, -16, -43, 4, -17, 4, 51, 23, -7, 1, -6, -48, -53, -35, -15, 4, 19, 12, -30, 38, 16, -6, 13, 5, -12, 23, -2, 0, -56, -71, -47, 14, 1, 42, 41, 4, -26, -1, -29, -72, -90, -51, -42, 4, 49, 46, 19, 45, 8, 3, 0, -37, -2, 38, 34, 31, -39, -48, -43, 6, 21, 59, 57, 0, -15, -42, -46, -74, -37, -38, -38, 34, 59, 64, 54, 65, 11, -30, -37, -41, -30, 19, 27, -8, -4, 13, -27, -24, -2, 57, 58, 2, -21, -32, -33, -54, -45, -30, 8, 66, 50, 40, 60, 68, 16, -14, -10, -48, -48, -43, -5, -15, 34, -4, -16, -32, 16, 63, 57, 8, -53, -42, 0, -26, -1, 11, 23, 31, 50, 83, 68, 45, 0, -29, -38, -41, -64, -59, -54, -27, -44, -22, -58, -47, -1, 47, 81, 21, -78, -43, -5, 22, 33, 18, 43, 19, 11, 13, 65, 103, 54, 25, -37, -17, -44, -28, -27, -60, -43, 23, -28, -19, -26, 39, 104, 42, -1, -13, 7, 28, 52, 49, 32, 32, 47, 41, 93, 105, 52, -4, -40, -11, -19, -58, -44, -29, -17, 34, -46, -5, -13, 54, -6, 19, 22, 32, 24, 59, 8, 76, 11, 8, 10, 54, 146, 102, 27, -67, -79, -48, -29, -4, -26, 6, 34, 29, -46, -15, 0, 48, 7, -39, 21, 36, 55, 51, 63, 23, -19, -35, -35, 95, 149, 122, 19, -102, -90, -39, -35, 24, -12, 29, 20, 37, 22, -20, -35, 2, -56, -138, -44, 40, 20, -20, 41, 13, 0, -20, -3, 89, 188, 104, -25, -106, -85, -79, -10, 35, 30, 31, 15, -3, -47, -50, -11, -36, -6, -73, -67, 0, 27, -22, 18, 40, 5, 9, 18, 97, 131, 59, -40, -100, -60, -31, 18, 45, 8, 8, 9, 9, -26, -23, -10, 24, 33, -84, -75, -64, -10, -15, -29, 5, -23, -19, 15, 69, 87, 41, -36, -67, -37, -38, -15, -7, -19, -37, 60, 37, -30, -15, -33, 15, 11, -27, -35, -58, -18, -17, -19, -51, -36, -37, 36, 75, 62, 30, -42, -60, -60, -33, -2, -73, -63, -88, 39, 56, 36, 3, 19, 6, 4, -50, -29, -9, -19, -30, -23, -15, -19, 24, 56, 114, 65, 57, -3, -16, -7, -40, -31, -79, -49, -88, 19, 67, 17, -18, -13, -23, 38, 20, -23, -39, -35, -25, 15, 21, -13, 3, 52, 59, 73, 10, 16, -29, -67, -67, -61, -45, -4, 9, 43, -17, 45, 3, -20, 15, -4, -24, -67, -60, -58, -31, -36, 22, 4, 21, -16, 3, 36, -10, -18, -22, -27, -12, 29, -6, 27, 44, -26, -1, 3, 16, -7, -18, -34, 1, 10, 30, -1, -9, 2, 39, 46, 29, 14, 42, -8, -26, -20, -27, -18, -15, -42, 33, 68, 20, -36, 2, -1, 16, -17, 2, -21, 39, 22, -17, -18, -11, 4, -13, 43, -10, -36, -18, -27, -48, -25, -24, -15, 14, 19, 29, 54, 13, -3, 15, -11, -6, 3, -3, -6, -12, -19, -8, 24, -9, 4, 32, 20, 5, 17, -38, -61, -71, -41, -31, -24, -7, 3, 27, 58, -16, -18, -5, 2, 13, 20, 14, -9, -6, 13, 2, -3, -16, 19, -19, 20, 18, -12, 13, 31, -18, 11, -11, 14, -18, 1, -19, -2, 8, -9, 1, -10, 15, 10, -441, 14, -13, 20, 3, -37, -8, -35, 4, -14, -37, -59, -8, 17, -25, -92, -19, -23, -54, -38, -23, 6, -15, -44, -23, 14, -13, 13, -5, 10, -14, 16, 13, 30, 9, -16, 20, -64, -9, 15, -6, -21, -14, -21, -10, 2, -3, 6, 15, 28, 70, 47, 56, 6, -15, -9, 5, 11, -29, 13, -23, 7, -3, 3, -5, -34, -55, -72, -51, -53, -24, -61, -55, -25, -26, -41, -19, -45, -12, -1, -51, -30, 21, 11, -9, -15, -20, -25, -34, 25, 18, 18, 3, -4, -35, -63, -19, -54, -56, -11, -30, 16, 34, 9, -34, -35, -65, -33, -40, -46, -45, -2, 19, -17, -8, -26, -38, 2, 24, 45, 9, 9, -5, -1, 2, 6, 0, 34, 1, -10, 24, -1, 11, -41, -19, -12, -57, -10, -53, -2, 12, 4, -21, -32, -27, -29, -40, 13, -6, 5, 6, -41, -1, -6, 5, 3, -24, -26, 1, -35, -20, -3, 28, 25, 4, -37, -27, -1, 22, -12, -28, -23, -59, -59, -52, -43, 2, -31, -20, -13, 1, -23, -50, -57, -32, -49, -40, -44, -60, -30, -6, 19, -2, -6, 14, 16, 16, -18, -2, -33, -91, -100, -49, -25, -18, -6, 14, 28, -1, -31, -37, -60, -54, -43, -52, -80, -75, -43, -54, -21, -13, -46, -20, -10, -20, -8, -12, -40, -112, -119, -51, -51, -36, -9, -2, -21, -44, -41, -21, -47, -32, -46, -15, -47, -43, -52, -71, -17, -32, -37, -51, -33, -1, -28, -7, -74, -99, -107, -81, -48, -31, -35, -26, -38, -54, -43, -13, 17, 24, 27, 2, 46, -3, -51, -81, -112, -74, -25, 22, -4, 3, -46, -41, -71, -65, -79, -111, -63, -52, -39, -7, 1, -6, -2, 51, 46, 52, 52, 66, 66, 63, -2, -100, -102, -55, -17, 35, 30, -4, -48, -55, -50, -66, -67, -117, -86, -36, -10, 16, 18, 23, 19, 21, 18, 38, 60, 11, 37, 94, 21, -52, -102, -26, -25, -10, 31, 5, -29, -19, -13, -89, -86, -91, -115, -24, 50, 59, 45, 31, 4, 43, 41, 62, 52, 8, 7, 42, -2, -36, -64, 10, 1, -21, 39, 1, -13, -70, -54, -97, -174, -145, -86, 23, 90, 107, 65, 47, 25, 18, 76, 47, 8, -22, 5, -13, -20, -51, -47, 13, 0, -36, 12, -21, -25, -97, -64, -121, -145, -49, 36, 84, 119, 103, 64, 72, 78, 66, 84, 58, 37, 16, 42, 14, -27, -40, -22, 34, 16, 2, -20, -17, -34, -79, -99, -137, -93, -18, 52, 95, 126, 88, 73, 85, 100, 100, 143, 86, 54, 40, 17, 3, -9, 4, -31, 45, -7, -8, -30, -27, 18, -40, -102, -167, -120, -82, 9, 22, 38, 49, 55, 69, 62, 70, 57, 44, -16, -8, -13, -32, -40, -26, -28, -37, -16, -35, -37, -29, 19, -74, -94, -95, -102, -40, -11, -12, 3, 15, 3, 16, 27, 1, -47, -28, -29, -48, -46, -45, -77, -48, -82, -37, -17, -45, -47, -40, -19, -55, -16, -51, -77, -49, -16, -27, -14, -18, -24, 2, 1, -35, -52, -74, -58, -28, -58, -47, -36, -62, -60, -46, -10, -7, -58, -33, 17, 0, 17, -36, -67, -66, 11, -56, -16, -30, -46, -26, -42, -32, -21, -30, -29, -63, -38, -38, -42, -33, -40, -29, 11, 2, -61, 27, 14, 3, -13, -8, -10, -25, -16, -8, -49, -55, -56, -39, -27, -17, 3, -8, -49, -21, -12, -38, -20, -21, -45, 11, -14, -40, -68, 10, 15, -34, 1, -11, -12, -30, -50, -44, -44, -58, -17, 4, 15, -23, -17, 2, 18, 26, 17, 2, 55, -3, -1, -4, 1, -19, -1, 10, 32, -16, -6, 12, -18, -72, -53, -27, 18, -20, 5, -22, 39, 27, 23, 41, 39, 14, -21, -6, 65, 94, 88, 18, 13, 4, -19, 8, 21, -32, -61, -18, -43, -23, -26, -8, -1, -57, 4, 21, 7, -1, -9, -20, -27, -23, 1, 14, 9, 31, 73, 43, -35, -3, -2, -9, -21, -13, -8, -27, -41, -45, -48, -74, -70, -99, -46, -66, -74, -86, -105, -155, -118, -94, -91, -67, -90, -59, -8, -24, -33, -23, -8, 0, 4, -20, -33, -40, -32, 26, 37, -20, -68, -57, -65, -92, -97, -66, -71, -113, -82, -108, -92, -49, -55, -13, -17, -36, 1, -10, 20, -1, 13, 2, 8, -4, -23, -43, -7, -42, -38, 21, -82, -70, 3, 5, -26, -42, -37, -27, -20, -20, -37, -32, -23, -5, -6, 9, 2, -8, -13, -12, -14, 20, -13, -2, -16, 17, 9, -17, -14, 3, 11, 0, -3, -10, -8, -7, 20, -8, 10, 18, -15, -19, 8, -2, 19, 15, -620, 12, 3, -15, 1, -14, -22, -4, 18, -21, -3, 5, 4, 39, 37, -32, 5, -8, -8, -29, -6, 16, 14, -3, -19, -2, 5, -19, 5, 6, 18, 1, 13, 28, -16, 21, 21, -19, -22, -26, -55, -44, -68, -70, -35, -46, -98, -58, -86, 6, -8, 28, 39, -14, -6, -6, 7, -19, 34, 10, 20, 1, 35, 34, 10, -67, -79, -88, -127, -143, -133, -114, -104, -162, -160, -159, -141, -132, -101, -88, -50, -29, -23, -12, -21, 8, 51, 59, 51, -27, 29, 27, -10, -24, -22, -55, -93, -112, -151, -145, -130, -101, -96, -92, -116, -90, -40, -33, -98, -93, -17, 14, 17, 2, 29, 45, 42, 26, 53, 62, 56, 10, 2, -40, -9, -45, -48, -27, -25, -35, -29, 1, -56, -40, 35, 29, 36, -32, 7, 17, -1, -1, -8, 58, 70, 66, 54, 101, 94, 37, 52, 6, 6, -8, -21, -15, -2, -31, 14, 35, 15, 19, 21, 92, 112, 27, -35, 18, 0, 16, -6, 59, 97, 105, 63, 78, 65, 61, 66, 65, 18, -16, 21, 10, 17, 36, 29, 43, 9, 3, 16, 13, 48, -9, -41, -6, 0, 19, 87, 87, 95, 56, 77, 85, 69, 63, 71, 33, 24, 23, 29, -18, 40, 32, 37, -6, 38, 7, 14, -20, -2, 14, 38, -17, 12, 18, 66, 156, 32, 48, 26, 17, 70, 36, 7, -20, -20, -9, 16, 8, 32, 6, 18, 11, 28, 31, 18, -8, 16, 25, 19, -37, 15, 67, 5, 108, 27, 10, 28, 0, 30, -3, -13, -36, -28, 16, 53, 4, 25, -14, 32, 17, 29, 25, -1, -14, 32, 47, -25, -9, 9, 69, 50, 93, 7, 7, 6, -11, -37, -48, -17, -61, -21, 19, 41, 21, 35, 26, 55, 40, 0, 5, 8, -17, -18, 46, -35, -34, -1, 24, 90, 131, 21, -23, -13, 1, -54, -87, -50, -28, -2, 54, 84, 49, 47, 52, 42, 13, -36, 7, -13, -28, -44, 53, -35, -53, 5, 33, 48, 77, -20, -24, -40, -46, -57, -82, -51, -14, 22, 11, 50, 70, 10, 38, 6, -3, -14, -16, 7, -29, -34, 76, -39, -21, 26, 67, 105, 29, -33, -36, -41, -75, -80, -52, -24, -18, 2, 21, 11, 8, -2, -26, -2, -31, -24, -14, -11, -68, 18, 93, -38, -64, 30, 70, 84, 14, -21, -37, -34, -7, -42, -23, -20, -23, -24, -15, 25, 9, -15, -25, -26, -37, -19, -27, 9, -13, -7, 39, -13, -22, 11, 48, 17, 51, -42, -41, -27, -10, -39, -46, -22, -31, -27, -52, -17, -32, -36, -23, -23, -39, -18, 22, 46, 25, 10, -30, -22, -33, 16, -21, -13, 43, -55, -59, -71, -36, -41, -30, -80, -86, -35, -39, -24, -29, -23, -11, -21, -24, -16, 24, 12, 34, -25, -78, -8, -14, -27, -18, 8, 17, -39, -74, -53, -38, -42, -55, -86, -73, -51, -18, 13, -7, 15, 29, 0, -39, -22, 3, -15, -6, -54, -81, -45, -33, -33, -16, -4, -27, -31, -37, -50, -42, -56, -92, -83, -75, -56, -32, -26, 20, 21, 31, 18, -24, -31, -57, -85, -72, -89, -56, -40, -45, 5, 0, -16, -54, -5, -22, -28, -56, -48, -30, -59, -12, -41, -23, 9, 4, 7, 30, 23, -15, -42, -64, -53, -127, -92, -86, -7, 25, -20, 17, -32, 31, 1, -45, 27, 15, 5, -6, -28, -31, -29, -27, -12, -19, 7, 14, -25, -56, -64, -52, -89, -121, -116, -73, -46, -57, -12, 34, -16, 48, 14, 8, 3, 22, 18, 10, 27, -17, -8, 3, -9, -47, -34, -29, -10, -51, -72, -75, -71, -114, -47, -62, -27, 4, 5, 20, 6, 40, 74, 17, 32, 57, 41, 56, 57, 4, -16, -4, -7, -17, -21, -30, -25, -48, -43, -81, -52, -13, 2, -23, 46, -7, 12, 6, -22, -29, -16, 38, 6, 8, 25, 8, 2, 7, 26, -2, 3, -34, -26, -82, -33, -54, -23, -55, -35, -45, 9, -47, 2, -20, 14, 16, 8, 9, 51, 41, 58, 22, -42, 6, -9, -20, -15, -29, -62, -16, -45, -57, -46, 18, -33, -24, -19, -40, 12, -6, 11, -13, 1, -14, 10, 31, 71, 78, 68, 79, 81, 68, 43, 39, 38, 80, 43, 67, 74, 83, 117, 120, 101, 46, 47, 16, 20, 1, 9, -4, -5, 8, 11, -5, 12, 51, 33, 48, 75, 35, 88, 46, 53, 78, 15, 18, 68, 57, 57, 49, 42, 41, 31, 16, 11, -2, -19, -13, 19, 1, 19, -4, -12, 18, -8, -17, 7, 19, -1, 5, 7, 19, 9, 30, 14, 2, -9, 2, -1, -7, 1, -16, -2, 8, -7, 2, 13, 103, 18, -13, -5, 4, 23, 14, 33, 1, -21, -14, -16, -1, -26, -28, 35, -22, -20, 38, -11, -7, 3, -26, 15, 14, -13, 6, 15, 11, 1, -20, 3, -12, -6, 10, 9, 2, 30, 9, -13, -3, 12, -5, 12, 5, 6, -1, -12, 1, -22, -69, -81, -98, -4, -12, -8, -3, 8, 12, 11, -67, -83, -56, -14, -12, 14, 11, 4, 73, 46, 46, 50, 43, 25, 38, 16, 41, 14, 22, -16, 18, -24, 8, -17, 12, 0, 17, 9, -20, -76, -33, -14, 15, 15, 13, 31, 90, 81, 64, 47, 55, 22, 14, -15, 7, -13, -16, -45, 5, 46, 16, -11, -7, -7, -32, -34, -31, -6, 29, 15, -13, -33, 2, 27, 75, 70, 28, 40, -3, 20, -55, -28, -47, 15, -4, -54, 37, 39, 61, 0, -13, 3, -13, -7, -36, -19, 58, 15, -39, 17, -4, 18, 27, 77, 30, 37, -6, 12, -6, -22, -17, -1, 21, 24, 29, 43, 74, -10, -11, -13, 8, -16, -47, -6, 75, 27, 3, 41, -7, 45, 57, 27, 25, 32, 4, 19, -2, 27, 18, 21, 60, 36, 70, 56, 65, 8, -7, -1, -13, -16, -4, 4, 14, 53, 35, 24, 42, 8, 17, 33, -13, -5, -13, 43, 44, 36, 36, 39, 22, 48, 81, 67, 23, -3, 5, -24, -27, -11, 15, 48, 76, 56, 86, 63, 65, 72, 13, -2, -34, -44, 1, 37, 77, 38, 40, 13, 36, 61, 71, 102, 33, 4, -15, -21, -10, 17, 73, 64, 66, 89, 102, 114, 117, 38, 12, -27, -53, -46, 9, 10, 7, 10, 33, 0, 0, 21, 39, 102, 35, 5, 2, 50, 22, 36, 63, 67, 23, 55, 68, 98, 69, -2, -15, -64, -36, -41, -14, 4, -4, 4, 20, 22, -1, 4, 30, 48, 53, 0, -9, 49, 81, 85, 70, 54, 49, 21, 61, 31, 36, -22, -30, -42, -52, -34, -1, -18, 1, 12, 13, 36, 35, 5, 13, 39, 55, 5, 25, 33, 42, 90, 59, 36, 23, 51, 68, 74, 12, 1, -4, -27, -27, -6, -14, 6, -48, -18, -3, 48, 58, 50, 30, 34, 35, -6, 5, 44, 98, 49, 80, 86, 93, 82, 62, 74, 19, 20, -18, -8, -17, -34, -56, -29, -44, -74, -35, -2, 73, 73, 75, 33, 49, -18, -37, 26, 95, 73, 103, 142, 91, 79, 81, 84, 56, 32, 29, -1, -54, -98, -93, -20, -51, -19, -58, -59, 48, 94, 46, 82, 63, 29, -14, 56, 22, 31, 75, 70, 84, 59, 56, 69, 28, 20, 7, -44, -77, -105, -63, -42, -21, -15, -30, -12, 68, 120, 81, 83, 35, 41, 8, 36, 3, -52, -41, -18, 8, 4, 36, 21, 11, 24, -13, -23, -24, -56, -50, 2, 15, 24, -8, 48, 96, 105, 74, 72, 52, 23, 28, -5, -13, -124, -73, 0, 11, -9, -5, -34, 4, -2, -8, -56, -19, -34, -32, 38, 56, 52, 18, 73, 110, 46, 47, 73, 62, 11, 13, -15, 6, -10, -56, 16, 11, 26, -5, -14, -23, -20, -11, -58, -58, -50, 3, 35, 43, 42, 13, 74, 73, 42, 47, 73, 62, 39, 29, 42, 32, -71, -49, -5, 15, -16, -21, -39, -23, -11, -20, -18, -45, -14, 10, 49, 51, 23, 3, 7, 30, 0, 14, 42, 57, 56, 16, 31, 4, -35, -21, -43, -23, -16, -34, -36, -26, -46, -41, -23, -28, -8, 8, 49, 17, 27, 37, 62, 68, 0, -8, 7, 35, 81, 14, 8, -23, -6, -65, -66, -31, -15, -19, 12, -4, 31, 33, 40, 4, 22, 21, 59, 27, 50, 84, 93, 58, -1, -3, -1, 26, 28, 17, 25, 49, 41, -25, -20, -14, 51, 26, 53, 66, 90, 90, 29, 33, 64, 78, 66, 92, 70, 81, 10, 6, -42, -24, -28, -21, -11, -14, 45, 52, 42, 17, -22, 15, 56, 100, 62, 56, 78, 81, 74, 89, 45, 104, 99, 105, 60, 37, 25, 6, -14, -34, -13, -11, 10, -20, -1, 4, -6, 88, 98, 101, 88, 129, 93, 117, 112, 161, 136, 142, 169, 95, 129, 114, 68, 78, 37, 49, 33, 21, -9, -16, -16, -4, -2, 7, 29, 59, 57, 65, 85, 46, 35, 92, 92, 134, 93, 117, 70, 64, 101, 89, 65, 54, 4, 29, 17, 9, 28, 20, -14, -14, -18, 15, 4, 3, -2, 32, 21, 60, 32, 38, 59, 78, 17, 21, 44, 7, 19, 28, 18, 0, 27, 0, 21, 10, -19, 7, 20, 11, 0, 13, 9, -8, -19, 3, 16, -11, -4, -13, -7, 19, -3, 0, 22, 17, -3, 18, -17, 8, -1, -6, 19, -12, 8, -20, 3, -9, -1280, 11, -17, -6, -12, -22, -25, -38, -3, 30, 41, -10, 19, 20, 28, -23, -28, 9, 19, 15, -18, -3, -16, -33, -11, 13, 18, 15, -16, -14, 8, -21, -20, -16, -68, -42, -21, -22, -12, 28, 14, 7, -22, -59, -4, 6, -7, 12, -12, -13, 12, 39, 51, 11, -17, -15, -1, 19, -20, -24, -22, -16, -6, -63, -36, -92, -48, -5, -49, -55, -22, -55, -87, -93, -76, -38, -22, -30, -53, -64, -37, -22, -17, 11, 2, -17, 22, 46, 18, 55, 23, -4, -13, 3, 12, -9, -48, -48, -60, -69, -68, -25, -21, -60, -62, -9, 4, 17, -55, -61, -51, 19, 16, 15, 53, 8, 27, -32, -13, 14, 47, 42, 76, 86, -1, -15, -48, -35, -2, -63, -21, -58, -23, -36, 16, 40, -59, -48, -50, 17, -5, 9, 43, 5, 21, 7, -18, 51, 70, 73, 99, 61, 21, -10, 6, -32, -43, -88, -29, -17, -3, 0, 11, 74, -6, -28, -24, 19, 10, 4, 5, 40, 81, 49, 17, 90, 54, 82, 101, 34, 35, -10, -22, -28, -23, -7, 10, -11, 12, -1, -18, 12, -47, -74, -46, 8, 3, 22, 49, 102, 89, 86, 89, 84, 67, 69, 71, 47, 49, -37, -6, -41, 3, 29, 8, -10, 13, -11, -11, -92, -70, -89, -58, -41, 19, 58, 60, 88, 81, 124, 83, 64, 44, 25, -9, -31, -1, -56, -6, 22, 10, 26, 21, 58, 3, 4, -57, -105, -94, -35, -48, -34, 18, 44, -9, 41, 48, 76, 93, 54, 5, -31, -88, -84, -87, -43, 20, -8, -4, 32, 34, 71, 37, -66, -154, -137, -62, -18, -54, 22, -43, -10, -7, 26, 39, 37, -10, -3, -63, -140, -138, -126, -59, -30, 19, 5, 10, 0, 57, 26, 9, -91, -140, -129, -53, -56, -30, 21, 12, 16, 7, -23, 9, 15, -9, -36, -115, -190, -165, -84, 13, -12, 8, -28, 16, 59, 53, 22, 8, -72, -138, -127, -40, -30, 22, 19, -13, 50, 77, -21, -28, 25, -31, -74, -184, -211, -148, 6, 52, 2, -4, 28, -2, 22, 8, -16, -8, -121, -161, -131, -37, -45, 0, -17, -6, 32, 45, 15, -18, -37, -48, -107, -174, -161, 19, 60, 72, 45, 5, 13, -4, -19, -1, 13, -23, -79, -162, -137, -49, -11, -34, -20, -18, 38, -46, -37, -79, -74, -86, -114, -159, -91, 85, 116, 101, 60, 15, 53, 0, -19, 19, -13, -1, -43, -100, -56, -26, -35, -43, -31, 15, -15, -71, -60, -115, -111, -172, -146, -141, -18, 100, 87, 88, 90, 64, 32, 46, 58, 32, 30, -37, -68, -57, -85, -61, -103, -1, -16, -7, -23, -70, -137, -202, -181, -193, -99, -96, 23, 49, 60, 65, 74, 59, 35, 78, 79, 45, 1, -44, -50, -74, -112, -101, -105, 7, -14, -23, -16, -39, -142, -115, -123, -114, -78, -84, -36, -22, 0, 38, 99, 45, 22, 59, 57, 10, -61, -49, -81, -150, -108, -122, -91, -48, 1, -31, -1, -104, -111, -55, -56, -17, -52, -70, -66, -50, -50, 5, 20, -10, 21, -6, 36, 5, -43, -44, -81, -114, -99, -76, -62, -26, -67, -37, -65, -95, -45, -83, -70, -10, -60, -79, -43, -75, -23, -15, 18, -14, -1, 4, -6, -37, -78, -65, -67, -51, -86, -83, -94, -69, -57, -23, 8, -42, -78, -73, 7, -6, -25, 4, -3, -22, 1, -14, -5, 20, -9, -23, -14, -42, -58, -75, -87, -118, -115, -101, -107, -57, -63, -3, -1, -44, -85, -15, -11, 19, -5, -50, -35, 8, -7, -22, -28, -16, -44, -48, -55, -77, -69, -67, -87, -67, -82, -73, -45, -73, -28, 10, -14, -31, -90, -19, 1, 11, 15, -37, -22, -29, -49, -8, 14, 9, -14, -69, -71, -65, -130, -71, -1, 23, 12, 16, -31, 34, -2, -6, -42, -75, -111, -98, -66, -23, -1, -18, 21, -28, -7, 31, 30, -1, -7, -37, -79, -48, -46, -32, -21, -9, -11, -1, -22, 9, -20, 1, -14, -49, -51, -28, -60, -49, -47, -127, -82, -50, -10, 18, 36, 24, -17, -86, -58, -61, -47, -84, -61, -64, -57, 7, 32, 34, -17, 13, -12, 12, 10, -1, -16, 10, 22, -26, -68, -50, 38, 76, 91, 79, 35, 41, -27, -7, 32, 23, 8, 26, 20, 12, -17, -19, -16, -9, -2, -9, -11, -3, -27, -19, -20, -41, -27, 6, -42, -20, 13, 25, -53, -31, -3, -14, 9, -22, -21, -20, 4, 18, -2, 2, -11, 14, -15, -3, 13, 8, 16, -3, 13, 19, 11, -20, -19, 8, 1, -3, -7, 7, -1, 14, -8, 12, -5, -7, -5, -2, -7, -18, 12, -9, 792, 6, -19, -17, 8, -25, -1, -35, 1, -14, -29, -49, -5, 33, 8, -48, 15, 2, -68, -43, -30, 6, 16, -13, 7, -11, 7, 6, 11, 16, -13, -19, 27, 9, -9, -21, -8, -65, -12, -5, 8, 9, 25, 8, 31, 5, -1, 48, 50, 32, 41, 62, 91, 3, 0, 15, -17, -9, -9, -11, 22, 64, 38, 20, 37, 2, -34, -42, -15, -24, -16, 27, 33, 10, 28, 40, 65, 54, 38, 8, -19, -48, 55, -17, -17, 10, 19, 43, 13, 122, 125, 49, 60, 20, 7, -20, -22, -67, -55, -54, -43, -1, 22, 27, 38, 29, 2, -13, 17, 41, 15, 16, -5, -5, 49, 41, 48, 125, 111, 77, 123, 70, 20, 7, -6, -18, -41, -49, -60, -38, 25, 20, 10, -24, -14, 47, 47, 105, 68, 4, -9, -19, 3, 44, 59, 100, 60, 102, 91, 56, 43, 5, -23, -25, -44, -47, -19, -3, 10, 12, -23, -22, -35, -11, 98, 95, 24, -8, 9, 6, -52, 17, 48, 88, 57, 77, 62, 43, 59, 27, 17, -4, -6, -18, -33, -18, 1, 5, -16, 2, -46, -14, 48, 68, -3, 22, 12, -10, 12, 45, 48, 70, 50, 56, 75, 74, 81, 55, 66, 21, 14, -24, -62, -49, -28, -5, -32, -29, 28, 1, 15, 50, -6, -18, -3, -32, -9, 4, 28, 4, 9, 36, 2, 62, 69, 54, 69, 45, -7, -26, -55, -34, -6, -21, -5, -17, 24, 23, 6, 73, -53, -25, -11, -13, -56, 8, 5, -19, -17, 30, 32, 76, 50, 44, 34, 28, 0, 1, -18, -70, -63, -30, -34, 20, 16, 5, 26, 131, 10, 24, -36, -63, -61, -10, -62, -38, -8, -3, 42, 75, 46, 10, 44, 41, 31, -1, -37, -58, -42, -54, -22, 29, 14, 32, 27, 95, 23, 39, -12, -42, -50, 22, 1, -44, 8, -25, -25, 17, 46, -11, 59, 30, 77, 80, 10, 3, -32, -4, 0, 19, 44, 60, 25, 75, 9, 33, 8, -22, -41, 1, -75, -70, -23, -36, -49, -12, 9, 44, 103, 87, 118, 94, 65, 5, 3, -5, 31, 12, 55, 49, 64, 69, -16, 7, -26, -31, -67, -13, -61, -32, -9, -15, -1, 8, -13, 41, 113, 104, 105, 108, 71, 6, -21, 26, 48, 18, 69, 25, 103, 101, -64, 7, 5, -35, -40, -47, -17, -27, -17, 0, 28, 44, 16, 30, 71, 92, 155, 140, 68, 19, 27, 58, 38, 65, 47, 53, 66, 92, -73, -33, 16, -30, -48, -64, -5, 8, -37, -6, 18, 36, 27, 36, 31, 63, 107, 84, 21, 21, 31, 21, 27, 49, 48, 64, 60, 49, -29, -24, -9, -1, -101, -80, -10, -16, -31, -32, 0, 18, 11, 15, -8, 11, -10, -33, -32, -35, -21, 11, 29, 10, 42, 63, 71, -14, -25, -54, -19, -68, -90, -43, -38, -39, -20, -29, -10, 13, -32, -56, -56, -70, -117, -101, -60, -45, -39, -42, 21, 24, -6, 8, 7, -29, -91, -52, -46, -32, -57, -57, -20, -38, -9, -6, -27, -26, -32, -78, -65, -57, -86, -52, -58, -40, -35, -48, -25, -26, -9, -42, -21, -24, -52, -35, -36, -42, 7, 56, -4, -62, -22, -26, -47, -24, -63, -28, -8, -35, -33, -45, -42, -36, -58, -49, -69, -36, -33, -34, -6, -2, -69, -60, -36, 23, 30, 46, -22, -36, -34, -21, -40, -43, -70, -30, -19, 7, 10, -43, -52, -37, -74, -41, -22, -25, -80, -13, 21, -37, -77, -40, -13, 38, 33, 84, 73, 21, -17, -60, 20, -20, -27, -18, -13, 19, -6, -56, -35, -39, -25, -25, -54, -47, -57, -87, 9, -33, -11, -6, 13, 38, 0, 9, 65, 92, 17, 25, 66, 42, 41, 32, 50, 25, -4, -16, 21, 10, 30, 4, -24, 0, 20, 11, 76, -1, 7, 15, 1, -4, -53, 1, 62, 34, 16, 35, 48, 71, 72, 45, 38, 49, 66, 73, 70, 55, 37, 29, 81, 101, 111, 73, 15, -27, 5, -14, 13, -8, 16, -40, 9, 22, -6, 29, 10, 39, 38, -6, 7, 24, 51, 33, 41, 18, 53, 27, 59, 65, 79, 20, 15, -27, 9, 8, 17, 10, -1, -46, -20, 5, 82, 83, 102, 78, 33, 65, 25, 78, 128, 96, 78, 97, 58, 53, 24, -1, 18, 10, 4, -22, -2, -1, 17, 7, 2, -1, 8, 10, 32, 33, 51, 15, 46, -20, -40, -26, 61, 13, -8, -4, 36, 24, -7, 11, 2, 22, 6, -2, -15, -3, 19, -12, -19, -16, 8, 19, 19, 15, -13, 3, -15, 0, 2, 19, 3, -18, -4, -19, 7, 14, -1, -17, -6, -12, 20, 7, -14, -2, 14};
    localparam integer positions[0:784][1:3] = '{
'{0,100480,108736},
'{785,100609,108801},
'{1570,100738,108866},
'{2355,100867,108931},
'{3140,100996,108996},
'{3925,101125,109061},
'{4710,101254,109126},
'{5495,101383,109191},
'{6280,101512,109256},
'{7065,101641,109321},
'{7850,101770,109386},
'{8635,101899,0},
'{9420,102028,0},
'{10205,102157,0},
'{10990,102286,0},
'{11775,102415,0},
'{12560,102544,0},
'{13345,102673,0},
'{14130,102802,0},
'{14915,102931,0},
'{15700,103060,0},
'{16485,103189,0},
'{17270,103318,0},
'{18055,103447,0},
'{18840,103576,0},
'{19625,103705,0},
'{20410,103834,0},
'{21195,103963,0},
'{21980,104092,0},
'{22765,104221,0},
'{23550,104350,0},
'{24335,104479,0},
'{25120,104608,0},
'{25905,104737,0},
'{26690,104866,0},
'{27475,104995,0},
'{28260,105124,0},
'{29045,105253,0},
'{29830,105382,0},
'{30615,105511,0},
'{31400,105640,0},
'{32185,105769,0},
'{32970,105898,0},
'{33755,106027,0},
'{34540,106156,0},
'{35325,106285,0},
'{36110,106414,0},
'{36895,106543,0},
'{37680,106672,0},
'{38465,106801,0},
'{39250,106930,0},
'{40035,107059,0},
'{40820,107188,0},
'{41605,107317,0},
'{42390,107446,0},
'{43175,107575,0},
'{43960,107704,0},
'{44745,107833,0},
'{45530,107962,0},
'{46315,108091,0},
'{47100,108220,0},
'{47885,108349,0},
'{48670,108478,0},
'{49455,108607,0},
'{50240,108736,0},
'{51025,0,0},
'{51810,0,0},
'{52595,0,0},
'{53380,0,0},
'{54165,0,0},
'{54950,0,0},
'{55735,0,0},
'{56520,0,0},
'{57305,0,0},
'{58090,0,0},
'{58875,0,0},
'{59660,0,0},
'{60445,0,0},
'{61230,0,0},
'{62015,0,0},
'{62800,0,0},
'{63585,0,0},
'{64370,0,0},
'{65155,0,0},
'{65940,0,0},
'{66725,0,0},
'{67510,0,0},
'{68295,0,0},
'{69080,0,0},
'{69865,0,0},
'{70650,0,0},
'{71435,0,0},
'{72220,0,0},
'{73005,0,0},
'{73790,0,0},
'{74575,0,0},
'{75360,0,0},
'{76145,0,0},
'{76930,0,0},
'{77715,0,0},
'{78500,0,0},
'{79285,0,0},
'{80070,0,0},
'{80855,0,0},
'{81640,0,0},
'{82425,0,0},
'{83210,0,0},
'{83995,0,0},
'{84780,0,0},
'{85565,0,0},
'{86350,0,0},
'{87135,0,0},
'{87920,0,0},
'{88705,0,0},
'{89490,0,0},
'{90275,0,0},
'{91060,0,0},
'{91845,0,0},
'{92630,0,0},
'{93415,0,0},
'{94200,0,0},
'{94985,0,0},
'{95770,0,0},
'{96555,0,0},
'{97340,0,0},
'{98125,0,0},
'{98910,0,0},
'{99695,0,0},
'{100480,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0},
'{0,0,0}
};

endpackage