package my_package;

    integer connection [89:0];

    localparam integer network_structure [2:0] = '{4, 37, 49};  
    localparam integer connectionRange [3:0] = '{90,86,49,0};
    localparam integer weigths [2001:0] = '{1216, 105, 219, -46, -366, -418, -300, 173, 375, -376, 27, 39, 60, -65, -109, -332, 139, -247, 98, 200, 30, 139, -214, -37, 75, 99, 294, -117, -59, -129, 260, -319, -410, -83, 48, -332, 263, 71, -483, 132, -35, 94, 348, -74, -126, 99, -362, 93, -12, -70, -116, -247, -151, 642, 286, -88, 80, -203, 201, -272, -188, 270, -299, 51, -215, -167, 94, 58, 21, 72, -25, 179, 34, -38, -264, 99, -1141, 49, -50, -240, -40, -408, 72, 90, -141, 311, -38, -39, -150, 249, 139, -524, -133, 285, -170, 4, 67, 0, 383, -222, 389, -60, -194, 62, 41, -143, -97, 64, 132, -6, 148, 221, 197, -267, 1827, -387, -323, 39, 217, 533, -66, -427, 214, 373, 81, 43, -17, 465, -69, 342, 222, 326, -151, -41, 218, 9, 133, 342, 72, -229, 244, -189, -311, -174, 249, -15, 210, -245, -382, 26, 114, 115, -7697, -2, 113, -2, 60, -55, -168, -181, 37, 113, 104, 5, -89, -85, -227, 115, 235, 261, 271, 134, -52, -139, 140, 171, 327, 354, 60, -57, -163, 183, 302, 314, 82, 94, 90, -94, -2, 165, 54, 32, 93, 88, -25, -133, -6, -13, -42, 87, -17, -58, -8468, -48, 124, -97, -10, 56, -43, -43, 38, 184, 4, -40, -122, -119, -80, 343, 170, 162, 23, -85, -62, 68, 119, 159, 32, -84, 41, -92, -87, 69, 136, 20, 131, 40, 28, -93, -147, 44, 117, -18, 69, 56, 122, -239, -152, -109, 225, 189, 32, -40, -4307, 91, 61, 88, 252, 144, 57, 278, 161, -54, -54, 171, -28, -169, 151, -53, -33, -76, -221, -51, -72, 2, -13, -184, 67, -90, 2, -14, 98, -87, -91, -56, -160, -138, -90, -55, 40, -9, 10, -12, -22, -79, -30, 81, 102, 128, 290, 151, 116, 31, 6032, 1, -150, 86, 77, 44, -144, -70, 48, -111, 168, 22, -27, 10, 28, -65, 38, -138, -192, 18, -75, -28, -56, -142, 4, -70, 79, 95, 41, 35, -247, -72, 62, -131, 81, 27, 210, -17, -78, -12, 36, -118, -29, 60, 45, 191, -33, 71, -38, -75, 8206, 6, -136, -224, -266, -177, -171, 9, -7, -131, -103, -468, -292, 45, -60, -25, -133, -84, -381, -167, -107, -115, 9, -29, -28, -158, -96, -127, -106, -171, -161, 10, 110, 68, -54, -15, -35, 11, 158, 173, 96, 20, 74, 208, 149, 140, 203, 101, 116, 148, -3465, -42, -80, 123, 46, 42, -82, -92, 70, 23, 61, 33, 101, 71, -118, -4, -29, -74, 108, -9, -102, -184, 101, 201, 69, 217, -42, -68, -118, 37, 139, 109, 108, 23, -81, -145, 41, 24, 54, 113, -122, -31, -274, 90, 103, 188, 26, 115, -108, -144, -7685, -114, -126, 8, -75, -72, -80, -196, -68, -41, -69, -73, -143, -152, -267, 55, 132, 82, 71, 159, 210, -32, 38, 8, 55, 363, 265, 129, -17, -9, 104, 187, 359, 297, 192, -19, -23, 198, 220, 261, 260, 239, 121, -65, -48, 37, 65, 247, 160, -3, 5401, 91, 75, -219, -255, -233, 28, 52, 114, -86, -248, -118, -21, -135, 53, 107, -114, -23, -32, -104, -16, 74, -71, 38, -29, -356, -270, -69, -25, 88, 161, -129, -237, -115, -143, -35, 182, 207, 154, 61, 60, 151, 180, 178, 159, -10, -15, -120, -24, 95, 12623, 139, -92, 142, -12, 20, -22, -88, -32, -63, 123, 151, 166, 170, -81, -204, -176, -140, -52, 26, -62, -165, 54, -35, -76, -59, -152, 0, -228, -67, -193, -73, 76, 82, -12, -107, 2, -54, 10, 29, 170, -12, -134, 227, 26, 145, -43, -61, -69, 42, 2346, 84, 131, 77, 80, 51, 54, 140, 132, 2, 87, 86, 90, 129, 59, 100, 60, 45, 65, 100, 73, 68, 77, 95, 71, 33, 86, 30, 34, 123, 50, 22, -10, -17, 34, 107, 116, 52, 27, 74, 93, 39, 101, 70, 131, 48, 59, 69, 44, 117, 2584, 104, 89, 17, 13, 61, 50, 57, 89, 124, 96, 90, 65, 61, 49, 87, 43, 120, 52, 108, 27, 74, 86, 20, 10, 16, 47, 5, 78, 38, 29, 102, 8, 56, 78, 48, 86, 116, 43, 15, 45, 14, 91, 89, 49, 121, 69, 106, 114, 67, -6676, -51, -53, -40, -18, -25, 141, 186, 49, -14, -173, -70, 13, 8, 95, 49, 90, 46, -39, -64, -74, 76, -110, 126, 283, 29, -29, -52, 109, -10, 141, 133, 121, 16, -174, 1, -16, -24, -65, -46, -77, -15, 140, -5, -38, -106, -28, -10, 120, 76, 10238, 120, 24, -45, -7, 28, 156, 174, 95, -4, 141, 258, 174, 81, 121, -1, -31, 46, 40, -102, -174, -111, 0, 20, 59, 70, -221, -91, -276, -217, 17, 203, 31, 56, -109, -162, -280, -219, 135, 151, -111, -42, -166, -208, -201, -75, -173, 5, -90, -12, -6574, -60, -58, 42, -46, -88, -79, -208, 33, 61, -36, -38, 64, 105, -136, -28, -129, 17, 106, -73, 12, -120, 162, 292, 94, 178, -18, -19, -73, 107, 196, 74, 38, 64, -1, -127, -42, 13, 115, 120, -9, 51, -110, 59, 29, 110, 1, 135, 46, -160, 6171, 71, 93, 66, 92, 70, -170, -106, 102, 23, 277, 169, -121, -251, -158, 147, 147, 108, -129, -95, -354, -227, 242, 102, -14, -291, 2, -74, 44, 190, 106, -152, -84, -329, 68, 142, 111, -90, -125, -48, 40, -198, -179, 36, -158, -4, 294, 67, -287, -197, 9079, 56, 42, -39, 8, -5, 59, 225, -29, -108, 73, 64, -94, -13, 30, 47, 65, -26, -183, 4, -40, 100, -51, -285, -42, -78, 2, -13, 71, -44, -289, -156, -62, -129, 11, 145, 111, -22, -163, -82, -1, 5, 115, 39, -50, -50, 51, 0, -19, 76, 10328, -3, -91, 89, -231, 4, -25, -15, -64, 73, -41, -147, 119, 143, 78, -50, -178, -166, 32, -139, 38, -62, 115, 14, -99, 144, -62, -79, -59, 1, 77, -13, 82, 41, -73, -57, 57, 82, 114, 186, -62, -22, -152, 121, 32, -3, -219, -68, -39, -69, -3131, -15, 94, -78, 43, -46, -55, -58, -33, 0, -41, 34, -107, -103, -21, 13, 102, 66, -106, 182, 44, 34, -66, -217, -8, -38, 133, 95, 207, 72, -118, -153, -4, 5, 39, 117, 41, 97, -90, -69, 198, -10, 86, 24, 50, -17, 63, 38, -63, -14, -4120, 42, 154, -16, -67, -96, 64, 135, -45, 104, -147, 69, 69, 85, -39, -28, -182, 156, 268, 144, 9, 1, -98, -94, 94, 151, 12, -27, -82, 50, 167, -68, -66, 35, -80, 52, 21, 151, -39, -156, -102, 75, 97, -7, 63, -96, -112, -130, 71, 43, 10523, 50, -54, -11, -86, -41, -129, -71, -108, -66, 154, 0, 23, 57, 13, -166, 18, -42, 8, -5, 76, -15, -89, -200, -197, -28, -18, 62, 72, -17, -246, -122, 12, -13, 144, 83, -34, -47, -72, -20, 31, 107, 121, 51, -24, -14, -149, 2, 107, 135, -2040, 65, 136, -41, -117, -62, 136, 28, 94, -5, -223, -38, 189, 64, 35, -17, -160, -15, 191, 122, 160, -5, -207, -85, 134, 152, 55, 58, -119, -7, 48, -29, 63, 154, -139, -108, 6, 82, 2, -78, -161, 68, 134, 5, 138, -19, -232, -110, 45, 72, 3396, -43, -96, 167, -115, 17, 44, -252, -99, 54, 64, -129, 114, 250, -101, -89, -130, -47, 45, -89, -5, -77, 149, 66, -94, 217, -109, -23, -204, 59, 70, 96, 158, 58, -37, -56, -7, 68, 51, 116, -66, 60, -65, -28, 26, 25, -187, -2, -54, -81, 10195, 102, -93, -80, -53, 20, 15, 181, -17, -19, -16, 4, -156, -108, 53, -61, -8, -12, -80, 27, -188, -46, 3, -201, 52, -54, 13, -45, 57, -76, -295, -49, 23, -17, -55, 99, 143, 17, -174, -49, -22, -17, 47, 132, 9, 41, 14, -16, -7, 177, 4733, -53, 32, -10, -254, -21, -9, -177, -79, 106, 45, -117, 187, 211, -73, -5, 25, 66, 197, 60, 70, 26, -22, 93, -171, -64, -198, -47, -164, 68, 110, 36, -66, 108, -59, -38, -87, 74, 178, 63, -55, 91, -79, -93, 42, 48, -262, -100, 45, -66, -4350, -18, 73, -53, 90, -57, -101, -48, -52, -72, 52, -19, -120, -96, -5, 19, 56, 3, 3, 215, 144, 97, -79, -159, -169, 4, 217, 81, 197, 8, -97, -116, -1, -39, 116, 59, 63, 125, -76, -116, 180, 104, 90, -29, 81, 49, 38, -100, 19, -34, 6357, 141, 103, -101, 1, -48, 131, 90, 110, -10, -250, -118, -94, -62, 5, 94, -3, -104, -219, -155, -53, 19, -89, -34, -117, -275, -273, -44, -22, 45, 43, -196, -239, -238, -98, 18, 59, 124, -45, -1, -63, -3, 188, 160, 134, 19, 63, 6, 119, 68, -6737, -126, -28, 103, -41, -40, -85, -92, -66, 121, -42, -24, 59, 96, -103, -34, -95, -5, 127, -38, 3, -16, 26, 162, -18, 216, 55, -5, -30, -18, 190, 91, 66, 120, -4, -49, -34, -57, 41, 165, 21, 89, -186, -113, 69, 72, 23, 40, 65, -38, -7560, 80, -88, 81, 39, -16, -150, -235, 108, -11, 63, -61, -114, -31, -189, 127, 82, 131, 41, 5, 41, -117, 112, 46, 231, 352, 60, 24, -8, 63, 8, 214, 82, 108, 193, 57, 73, -46, 45, -49, 11, 38, -112, -49, 7, -12, 12, 25, -13, -32, -5909, -9, -208, 87, 136, 16, -46, 29, 36, -93, 154, 135, -25, -78, -90, -34, -2, -4, 12, 57, -29, -104, 5, 14, 270, 320, 251, 47, 16, -54, -111, 117, 196, 95, 77, -40, -54, -137, -105, -4, -74, -164, -99, 66, -47, -45, 145, 86, -30, 19, 10665, 55, -10, -278, -286, -217, -6, 50, -34, -41, -116, -85, -47, -171, 90, 61, -26, -101, -172, -68, -206, 110, -46, -90, -94, -200, -234, -108, 4, 103, 13, -61, -95, -194, -64, 62, 174, 115, 101, 108, -3, 25, 58, 208, 226, 119, 156, -12, 70, 153, -1266, -13, -98, 185, 63, 183, -55, -8, -11, -41, 145, 28, 90, 136, -113, -50, -51, -57, 60, -80, -86, -146, 94, 112, 28, 130, -34, 30, -98, -2, -129, 36, 143, -64, -21, -65, 102, -65, -72, 32, -18, -124, -186, 234, 120, 173, -2, 24, -53, -131, 4411, -4, -99, 130, 32, 70, -21, 11, -88, -6, 90, -95, 109, 205, -33, -44, -52, -151, 22, -56, -125, -220, 141, 122, 29, 119, -138, -70, -162, -3, -18, 141, 111, 54, -71, -120, 55, 65, 29, 40, -60, -154, -169, 106, 91, 25, -62, -4, -43, -52, -5958, 40, -248, -62, 83, 4, -135, -91, 42, -36, 154, 31, 7, -19, -9, 73, 124, 77, 119, 88, -11, 36, 180, 90, 165, 285, 303, -18, 58, 138, -113, 154, 218, 123, 221, -5, 38, -88, -160, -81, 92, -55, -94, -45, -176, -131, -50, -37, -142, -115, -9166, -206, -156, 28, 22, 43, 59, -22, -116, -8, -19, -48, 96, 154, -85, -71, -14, 88, 197, 129, 352, 109, -157, -8, -52, 156, 307, 282, 71, -53, -41, 44, 140, 142, 191, 28, -134, 23, 173, 26, 144, 89, 24, -110, -53, 77, -3, 37, 116, -116, 1110, 16, -21, 190, -22, 154, 49, -146, -25, -18, 72, -63, 121, 225, -34, -53, -4, -125, 103, -76, -87, -142, 93, 140, -1, 183, -103, -95, -90, 19, -23, 24, 91, -21, -47, -50, 61, 43, 60, 50, -38, -150, -256, 54, 82, 111, -54, 10, -25, -150, 3550, -72, 128, -118, -144, -116, -19, -16, -1, 121, -105, -20, 128, 8, -46, 12, -38, 55, 43, 18, 137, 88, 1, 1, -114, -114, -180, -84, -68, 25, 185, 13, -145, 96, -82, -55, -30, 95, 188, 100, 0, 149, 93, -115, -11, -129, -235, -73, -33, 23, -1364, 117, -11, -45, 84, 110, 113, 348, 61, -6, -75, 104, -80, -109, 98, 98, -50, 48, -201, -116, -195, 122, -134, -46, 116, -167, 5, -124, 161, 7, 0, 81, -49, -143, 19, 51, 38, 28, 98, -13, -59, -136, 115, -2, -12, -32, 170, -6, 115, 89};

    localparam integer positions[0:49][1:2] = '{
        '{0,1850},
        '{50,1888},
        '{100,1926},
        '{150,1964},
        '{200,2002},
        '{250,0},
        '{300,0},
        '{350,0},
        '{400,0},
        '{450,0},
        '{500,0},
        '{550,0},
        '{600,0},
        '{650,0},
        '{700,0},
        '{750,0},
        '{800,0},
        '{850,0},
        '{900,0},
        '{950,0},
        '{1000,0},
        '{1050,0},
        '{1100,0},
        '{1150,0},
        '{1200,0},
        '{1250,0},
        '{1300,0},
        '{1350,0},
        '{1400,0},
        '{1450,0},
        '{1500,0},
        '{1550,0},
        '{1600,0},
        '{1650,0},
        '{1700,0},
        '{1750,0},
        '{1800,0},
        '{1850,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0}
    };

endpackage