package my_package;

    reg[31:0] connection [89:0];

    localparam integer network_structure [2:0] = '{4, 37, 49};  
    localparam integer connectionRange [3:0] = '{90,86,49,0};
    localparam [31:0] weigths [2001:0] = '{32'h3ca1867e, 32'hbf74a1a5, 32'h3dee22de, 32'h3ec23834, 32'hbe56fafe, 32'h3f11fd4a, 32'h3e085bc7, 32'hbf2b28bb, 32'h3f4ca6ac, 32'hbecc28b6, 32'h3f20f4d3, 32'h3eb60d93, 32'h3e7dc313, 32'h3f060b1c, 32'h3f18124e, 32'h3f355881, 32'hbf0aada5, 32'hbf7ef1c0, 32'hbf12abb3, 32'hbebd0777, 32'h3bcb76c0, 32'h3ebcd2b6, 32'h3ed6cb79, 32'hbf297ac3, 32'hbec26f3b, 32'h3e601f3d, 32'h3ece55fe, 32'h3dec2156, 32'h3f86cb8b, 32'hbf1ff41a, 32'h3f539485, 32'hbf4b6432, 32'hbf8c4989, 32'h3e392628, 32'h3e0de710, 32'hbf6669e8, 32'hbf33996a, 32'hbeb3c3c7, 32'hbc985974, 32'hbed1ef51, 32'hbf2732e4, 32'hbf17311f, 32'h3ec3906c, 32'h3ea85210, 32'h3edb01ad, 32'hbe2277bd, 32'hbebdea6f, 32'hbf05bfc7, 32'h3de08664, 32'hbebd9a71, 32'h3f4e8083, 32'hbf2942d0, 32'hbf49b695, 32'h3f27f33a, 32'hbe53ec5e, 32'h3f31c3f9, 32'hbd0d19c8, 32'hbe7fed47, 32'hbf5a6fdb, 32'h3e1a2ca5, 32'h3f456b2c, 32'h3eec750c, 32'h3d31918c, 32'hbf5c870a, 32'hbd4ae94e, 32'h3f9bb9ea, 32'hbecb5ead, 32'h3f818939, 32'hbf208b9b, 32'hbf3f2b56, 32'h3f94d5e3, 32'hbf68b022, 32'hbf4b1cfe, 32'h3f1f2dd2, 32'h3efdef56, 32'h3ecb532c, 32'hbd938207, 32'h3e66a304, 32'hbe95d8c5, 32'h3f48221c, 32'h3eb3a152, 32'hbf4f556d, 32'h3e9299b4, 32'h3f6a371d, 32'hbf924313, 32'hbdb75367, 32'hbebe6a36, 32'h3eee3a83, 32'hbe6afed4, 32'h3eba63f8, 32'hbd101564, 32'hbfaf15f3, 32'hbfdf8803, 32'h3f5d2a55, 32'hbd7e518d, 32'h3eb3d343, 32'h3f164b74, 32'h3e1f5b4f, 32'hbf2b1fb3, 32'hbf15d96c, 32'hbf0ed44b, 32'h3e546e36, 32'hbf394edd, 32'hbfad676a, 32'hbfb912a4, 32'hbfa44a30, 32'h3ed5effa, 32'h3f717600, 32'hbefd486e, 32'h3f22e88f, 32'h3f8a861b, 32'h3f42f5d0, 32'h3f1407f6, 32'h3d81cd37, 32'h3d26d179, 32'h3fa2742d, 32'hbf4efd8a, 32'h3f49d6be, 32'hbf45a9e5, 32'hbeaed3b1, 32'hbf8b6f88, 32'h3f219544, 32'h3fb98c0b, 32'h3fd582d0, 32'hbf3b203e, 32'h3e21c40d, 32'hbea737f1, 32'h3f1177a0, 32'hbec9efa8, 32'h3f50bef8, 32'h3fbc67f3, 32'h3f854b8d, 32'hbf207d0a, 32'hbf8b90cc, 32'hbf5e5857, 32'hbf37bbc9, 32'h3f4ac55a, 32'hbe9e571d, 32'h3ce09128, 32'hbf7a74c0, 32'hbeee9110, 32'h3f97c537, 32'h3f8d7440, 32'h3fbf925d, 32'h3f55affb, 32'h3fce6c28, 32'h3e7501f9, 32'h3f85354f, 32'h3eeb0c40, 32'h3f4a53b7, 32'h3e4e81ee, 32'hbf9e1b44, 32'h3f96641b, 32'h3e54330e, 32'hbe897e47, 32'hbee12718, 32'hbf47c09c, 32'hbe791d79, 32'h3d8f8ae2, 32'hbeb62a5b, 32'hbef4ee39, 32'hbe5df5e5, 32'h3e8ad334, 32'hbd162dea, 32'hbe153ecb, 32'h3ee6e144, 32'hbebe5e17, 32'hbe1ec165, 32'hbe311622, 32'h3f07c349, 32'h3d024754, 32'hbe9718e9, 32'hbefe0623, 32'hbe9f441f, 32'hbe5125ec, 32'h3ef23d5a, 32'h3f65a763, 32'h3f0532a7, 32'hbea49707, 32'hbf62cef4, 32'hbea414ec, 32'h3da071ae, 32'h3df65163, 32'h3ea043fc, 32'h3f0696e0, 32'h3eab0d84, 32'hbf15873a, 32'hbf43db21, 32'h3eb32fc9, 32'h3e20e112, 32'h3eafd56a, 32'h3e966a91, 32'hbe8d4814, 32'hbd2692dd, 32'hbee84957, 32'h3ee94017, 32'h3e9e7b29, 32'hbed81135, 32'hbf23b6b8, 32'hbf22350b, 32'hbf089550, 32'h3de65b31, 32'hbf8b645e, 32'hbda0ff36, 32'hbe877df2, 32'hbf0235a5, 32'hbe2cb606, 32'hbbe9d4ee, 32'h3d9b08a9, 32'h3e2faaa3, 32'h3d74dc5d, 32'hbde2ddee, 32'hbdb604e0, 32'hbe62b411, 32'h3f00ba24, 32'h3e2bd5c4, 32'hbddaf96c, 32'hbe2e356f, 32'h3db7057c, 32'h3f11dcc0, 32'h3e9f9cc8, 32'h3e383618, 32'h3e212d39, 32'h3f1cb915, 32'hbd2a7ffc, 32'h3eea691e, 32'h3e7b5141, 32'h3e4e7f61, 32'hbd890ee4, 32'hbe10c629, 32'h3d707f9e, 32'h3d6ca0c6, 32'h3f12d443, 32'h3eea42de, 32'hbea3994e, 32'h3ec9cd42, 32'hbe8bb521, 32'hbe821143, 32'hbd977033, 32'h3e6db108, 32'h3eccc9b1, 32'h3ea4761a, 32'hbdcf962c, 32'hbd546536, 32'hbcb51fe8, 32'hbe4f38f6, 32'hbe2aa9d1, 32'hbe102e2d, 32'h3e34152c, 32'h3e2ba88c, 32'hbe2bedf5, 32'hbdbbc958, 32'h3f19dac3, 32'hbe868c0a, 32'hbe026ff5, 32'hbec8edff, 32'hbef31e37, 32'hbde75408, 32'hbe383e84, 32'hbe6e5b1c, 32'hbf2b7838, 32'h3c44333f, 32'hbe62623f, 32'hbed8812b, 32'h3eb4eb50, 32'h3eedd9c7, 32'hbe4b29d7, 32'hbf045bb2, 32'hbcc945e1, 32'h3e94dbb8, 32'h3d83db87, 32'hbe791946, 32'h3cf48c19, 32'h3cf6c93d, 32'hbd883b75, 32'h3f0b139c, 32'hbedd6fe4, 32'hbeccf870, 32'hbec974ed, 32'h3b4115db, 32'hbe85692b, 32'hbea46650, 32'h3d825a29, 32'h3d97c6c5, 32'h3ca21412, 32'h3ec9d8fa, 32'h3dff0a15, 32'hbe015f1a, 32'h3d3f0b88, 32'h3f27531e, 32'h3f2fdc93, 32'h3ecca99b, 32'hbd965625, 32'h3e8827aa, 32'h3ef10def, 32'h3e2af84f, 32'hbca0d582, 32'hbe1a6633, 32'hbecbeeb9, 32'hbe90ae72, 32'hbe84fe36, 32'h3c88370c, 32'hbf1d7703, 32'h3e5650bb, 32'h3c804150, 32'h3f2d1db0, 32'h3ea91a0c, 32'hbdebf9a7, 32'hbe53acc6, 32'hbec2d8e1, 32'h3f0ac051, 32'h3f22fb71, 32'h3f04ae8b, 32'h3f05487c, 32'h3f291704, 32'h3e385b8c, 32'h3cd9e404, 32'h3f0c5a42, 32'h3eeb534a, 32'h3e3eca7f, 32'h3f4519d0, 32'h3e42307e, 32'h3d5c621d, 32'h3bcfa464, 32'h3f698c3f, 32'hbcd9ab3e, 32'h3f222cd1, 32'h3efc67a8, 32'h3f1068cf, 32'hbea39976, 32'h3e888ff9, 32'h3d8628e9, 32'hbe8fd733, 32'h3e0a32db, 32'h3f13a29c, 32'hbe918b86, 32'hbd9dc5b0, 32'hbe5cefbd, 32'h3e076540, 32'hbf0e12cf, 32'h3db39642, 32'hbdd9b5a9, 32'hbc598d0d, 32'hbeadc4ad, 32'hbef80fe5, 32'hbf0b6b44, 32'hbef0890b, 32'hbe568c0c, 32'hbe80a812, 32'hbeed357a, 32'hbeba7650, 32'hbeab0604, 32'hbd1d541a, 32'hbe8b6628, 32'hbd8421b6, 32'hbd81870e, 32'h3dd63486, 32'h3e9afbe7, 32'h3e8ea161, 32'h3e3c6a9a, 32'hbea0162d, 32'hbeca6e52, 32'hbdaf83a8, 32'hbe4fa595, 32'hbec4477b, 32'hbf424573, 32'h3e5062bf, 32'hbe5083f3, 32'h3e53bab0, 32'hbc1bfaeb, 32'hbe754af4, 32'h3f1f3573, 32'h3da411d5, 32'h3f083224, 32'hbf0c34f1, 32'hbee7141e, 32'hbe041ef8, 32'hbe828292, 32'h3e872755, 32'h3e564787, 32'hbd2e9820, 32'hbe58469a, 32'hbdea9f7e, 32'h3cd9d6d5, 32'h3c642632, 32'hbdb6ff87, 32'h3ecc4647, 32'h3eb3a632, 32'hbe0e76b8, 32'hbde11c47, 32'hbf33f26c, 32'hbf0dc6db, 32'h3e7762ef, 32'h3eb9db01, 32'h3ec7e904, 32'hbebd2b8c, 32'hbdf7b16a, 32'hbeca0b17, 32'hbe168cca, 32'h3eabce1c, 32'h3efb039d, 32'h3e889551, 32'hbf28e018, 32'hbb466995, 32'h3ee76203, 32'h3f473dec, 32'h3ea74b07, 32'hba131b70, 32'hbe68e8a4, 32'hbef2b12f, 32'h3ec47a72, 32'h3f3183f9, 32'h3f5c8cf2, 32'h3e161ad8, 32'h3ef2bb4d, 32'h3d86685b, 32'hbe314ee7, 32'h3f6bb3a0, 32'h3fb48182, 32'h3f76b9c7, 32'h3f8a65d8, 32'h3f0e3cfa, 32'hbe096801, 32'hbe4a592c, 32'h3ecab251, 32'h3ec21fb9, 32'h3faf3229, 32'h3f0a2198, 32'h3beef92e, 32'hbe9c76ca, 32'hbee05579, 32'h3daebe95, 32'h3dd78533, 32'h3ec427e1, 32'h3f09d034, 32'h3e1b38d3, 32'hbe447e7a, 32'hbe6d11cc, 32'hbe18b146, 32'h3e5f158a, 32'h3df0e4f0, 32'h3e5b5872, 32'h3df7dc66, 32'hbeaff56f, 32'hbefa1e7d, 32'hbec9aca3, 32'hbe1a9799, 32'hbb893dd7, 32'hbe2ceff2, 32'hbe817394, 32'hbf2b6f55, 32'hbf67af25, 32'h3f16aa2e, 32'hbe85e654, 32'h3cd91efe, 32'hba4c8735, 32'hbea84fa1, 32'hbe4f7e9b, 32'h3dc4ee39, 32'hbd123052, 32'hbee4a6bc, 32'hbc51c596, 32'h3edab76a, 32'h3e82a475, 32'h3af4a76d, 32'h3f04bd56, 32'hbea110f9, 32'hbed73375, 32'h3def41a8, 32'hbd90927e, 32'h3e4a543b, 32'hbe1f0f1e, 32'hbec2d36f, 32'hbee4f794, 32'h3ecc31c6, 32'h3edf54c1, 32'h3e7363f0, 32'hbe0c1ff8, 32'hbf1d91f8, 32'hbea81de5, 32'hbeb695b6, 32'hbedda277, 32'hbedb4ab7, 32'hbdcfd03a, 32'h3f01f7c5, 32'h3e5b71e9, 32'hbe232315, 32'hbe7db2d7, 32'h3e9149ee, 32'hbe11c189, 32'h3e7884dd, 32'h3f14ab5c, 32'hbdeebbdc, 32'h3e0c9a4b, 32'h3d5fa716, 32'h3df8df50, 32'hbbcfbba4, 32'hbdd820d6, 32'hbf05e1ff, 32'hbd7572e4, 32'hbe9cebe5, 32'h3c419a80, 32'h3f822d7b, 32'hbef98a47, 32'hbf02d42d, 32'hbf3e8f06, 32'hbeec3e3e, 32'hbf18c0c0, 32'h3ead723e, 32'h3e6bb662, 32'hbed85fea, 32'hbf6e3391, 32'hbf47be4d, 32'hbee23a64, 32'hbf0ebef9, 32'h3dde54b7, 32'h3d7afbbb, 32'hbf712572, 32'hbf411651, 32'hbe721d1c, 32'hbf72db60, 32'hbf1099e0, 32'h3d598edc, 32'hbde486db, 32'hbf4a6240, 32'hbea59830, 32'hbf3a2fb1, 32'hbf181fd6, 32'hbed8766a, 32'h3f1764ae, 32'h3d042718, 32'hbe989920, 32'h3e568c30, 32'h3e8ae6a2, 32'hbd84b0cd, 32'h3e6e3ba5, 32'hbcdd09a1, 32'h3f0d3d8e, 32'hbd5ef79b, 32'h3ebfe9ef, 32'hbdec5ff5, 32'h3e806e64, 32'h3eda9771, 32'h3ed16e6f, 32'h3f37d06c, 32'h3f25c7f3, 32'h3e95dc5b, 32'h3e16097c, 32'h3f34889f, 32'h3e77a513, 32'h3f22ff71, 32'h3f78388e, 32'h3f25176a, 32'h3e5a97d9, 32'hbe0f9c2b, 32'hbeec20da, 32'hbdc3005f, 32'h3e1ba153, 32'h3ee52316, 32'h3f1a218c, 32'hbed91880, 32'hbea81d1a, 32'hbeb501a2, 32'hbd74408d, 32'h3e900472, 32'h3eb54d3b, 32'h3f082189, 32'hbf1dbdb6, 32'hbf31d0d9, 32'hbf03a402, 32'hbf2145eb, 32'hbe2a1ee7, 32'h3ef4bc54, 32'h3ebe8076, 32'hbe9b432a, 32'hbf04a2b7, 32'hbf1eb417, 32'hbeac0a35, 32'hbdf5c379, 32'h3eae52b8, 32'h3df7a1e6, 32'hbf1d5eef, 32'hbeea3b91, 32'hbe676dc5, 32'hbd0bd1f4, 32'h3bfb5f80, 32'hbd891c00, 32'hbe17b391, 32'hbe101ff0, 32'hbf233253, 32'h3e250a73, 32'hbd14c1f7, 32'hbe7b0624, 32'hbd9d4c01, 32'h3dbbcddd, 32'h3cd621ce, 32'hbe37f630, 32'hbdd2e0dd, 32'hbd118f43, 32'hbeeb6ae4, 32'hbee4f8ce, 32'h3ebe8473, 32'hbf85910c, 32'hbee8e88b, 32'h3ebe8187, 32'hbcd13d1f, 32'h3f187d54, 32'h3dcd31dc, 32'hbebdd9b6, 32'hbe6c101c, 32'h3dca6263, 32'hbcc1277d, 32'h3dc87115, 32'hbe2ce5c9, 32'hbea2d48b, 32'hbeea1c6d, 32'h3e0d0439, 32'h3c62ce86, 32'h3eb3f596, 32'h3d9aa251, 32'h3e9ed3bd, 32'h3edc4aba, 32'h3f08610a, 32'h3e0ab98a, 32'hbebf3595, 32'hbcbb0ab6, 32'hbe856ece, 32'hbb76888f, 32'h3f58a7a0, 32'h3f05615d, 32'hbd57f843, 32'h3f2d41db, 32'h3d2e66d8, 32'hbd53e72e, 32'hbf6f4261, 32'hbe3af6b2, 32'h3e413902, 32'h3f06c2c6, 32'hbd87f712, 32'hbe2b2b02, 32'hbf15ae77, 32'hbed3d2f2, 32'hbc80c904, 32'h3d437b00, 32'h3f067b94, 32'hbe06e7e7, 32'hbcac7cf4, 32'h3e2935d7, 32'h3f1edd34, 32'h3ecc1127, 32'h3e55f9ca, 32'h3e845ea0, 32'h3f31825a, 32'h3da2ae9d, 32'h3e59dd48, 32'hbe084642, 32'hbf56e83c, 32'h3e5d52f5, 32'h3e57fa5e, 32'hbe08795c, 32'hbe35c93f, 32'h3e45b796, 32'hbdb20afa, 32'h3b51a3fe, 32'h3eb47084, 32'h3e7c3e71, 32'h3ccca95e, 32'hbe830d57, 32'hbde09ddd, 32'hbd7147a5, 32'hbca767ff, 32'h3e63f0b9, 32'h3f259bad, 32'h3ee9b741, 32'hbf202f0c, 32'h3e29bebe, 32'hbf656d18, 32'hbebd2223, 32'hbe661485, 32'h3e0f545c, 32'h3e809058, 32'hbf21ec6a, 32'hbe446336, 32'hbea2e823, 32'h3c3a3563, 32'h3f10d997, 32'h3dc0c65f, 32'h3dbc7648, 32'hbe4f1fee, 32'hbc0e0291, 32'hbd8d3287, 32'hbddc822b, 32'h3b2c172e, 32'h3ed45322, 32'h3e3252db, 32'hbe4db927, 32'hbdab086d, 32'hbe9079e8, 32'hbf6627ab, 32'hbd4397cc, 32'hbcbea1f2, 32'h3d9a7e4e, 32'h3e3d9ef8, 32'hbe80a3c7, 32'h3e69caff, 32'h3ea731a4, 32'h3d816e6c, 32'hbe83dcb5, 32'hbd319658, 32'h3e27e4bb, 32'h3e099f96, 32'hbe474748, 32'hbcb254af, 32'hbe15e598, 32'hbef02ca8, 32'hbe840e19, 32'h3d968772, 32'hbbfb74eb, 32'h3ece06b4, 32'hbe40231a, 32'hbe04abf1, 32'h3ed47f9d, 32'hbea9cf0b, 32'h3d3065e7, 32'hbe928381, 32'hbf365812, 32'h3d8b1d4a, 32'hbea4d1ac, 32'h3eb93bdb, 32'h3df32f9b, 32'h3d7574ab, 32'h3ea547cc, 32'hbec9b7e3, 32'hbed6b9c3, 32'h3da33889, 32'hbee316c0, 32'h3e93c37b, 32'h3e8ece97, 32'hbe2fe0dc, 32'hbdc843d4, 32'hbeea5f59, 32'hbe0f6a7b, 32'h3e270929, 32'h3ec6734d, 32'h3f1d7add, 32'hbeb4f9df, 32'hbef80e78, 32'h3e04a691, 32'hbe978c10, 32'h3e01317b, 32'h3ead6bba, 32'h3e536f95, 32'h3f03d9e7, 32'h3ddcfe43, 32'h3e0d6491, 32'h3e9c04ac, 32'hbe8ce8cc, 32'h3f03a161, 32'h3e8c5258, 32'h3e856761, 32'h3d94368e, 32'h3efbe055, 32'h3d20683b, 32'h3dc4ad92, 32'h3e461f3d, 32'h3f1df5e1, 32'h3f17c32f, 32'h3d7e4be2, 32'h3e09882b, 32'h3ed1149f, 32'h3bcf70f2, 32'hbe3ab680, 32'h3e8af6b6, 32'h3edb9142, 32'hbe9711d7, 32'hbdd0f9db, 32'hbf210a87, 32'hbf634814, 32'hbeaa189e, 32'hbe586856, 32'hbeeec60d, 32'hbecbfd03, 32'h3d5bc3f9, 32'h3a3813d9, 32'hbf59fe10, 32'h3f1beb25, 32'hbf1d52af, 32'hbe9eff72, 32'hbe8ff2b8, 32'h3eab55d5, 32'h3d0b83c5, 32'hbf2db657, 32'hbf3047f1, 32'hbf41c869, 32'h3d67db40, 32'hbe8ebd26, 32'h3c2388d8, 32'hbe6e2ead, 32'hbe739b23, 32'h3d487f87, 32'h3c3ec7df, 32'hbc9cec61, 32'hbf01a927, 32'hbdc392eb, 32'h3da5e153, 32'hbe097fa6, 32'h3d1b5e23, 32'h3e7ba3f3, 32'h3d31be6b, 32'h3ddec96e, 32'hbc03bc72, 32'hbd4c74d8, 32'hbe4f0349, 32'h3d995515, 32'h3f03dc39, 32'h3e25e8c0, 32'hbe9ccd1c, 32'hbe53beec, 32'hbd67ee1c, 32'h3f1b1a1a, 32'h3e9bbe1e, 32'hbd2af553, 32'h3f274191, 32'h3ecf44da, 32'hbe5eb5ca, 32'h3e7e2d55, 32'hbdaaf060, 32'h3db7c632, 32'hbd73e1a6, 32'hbde84c32, 32'hbe65f041, 32'h3dcc8aef, 32'h3f35ac9a, 32'h3f11b0f1, 32'hbef9c74d, 32'h3ee675f2, 32'hbe8187f3, 32'hbdbb5ccd, 32'hbe03ef0e, 32'h3e413250, 32'h3ee94e13, 32'hbeedc0ff, 32'h3d730eb8, 32'hbda0241f, 32'h3e9a8b7d, 32'hbdde7607, 32'hbd2bb60e, 32'hbef13200, 32'hbdd64deb, 32'hbdb15dc8, 32'hbbd6f542, 32'hbdd4bfcd, 32'h3edb5622, 32'h3f52a3d1, 32'h3f29678c, 32'h3e59b8c6, 32'h3f183c1a, 32'hbe85c921, 32'h3e7b5451, 32'h3e503a68, 32'h3f305590, 32'h3e5c4844, 32'hbe3c72e0, 32'hbe62dd2c, 32'hbf608bcc, 32'hbf837454, 32'hbe8baa45, 32'h3f155667, 32'h3c5266be, 32'h3d086b6f, 32'hbdcf335b, 32'h3eaae47c, 32'hbd060275, 32'hbd91a9b3, 32'h3e663cd4, 32'hbe1adf89, 32'h3ead43d6, 32'h3d50c13f, 32'h3da3e229, 32'hbe3f6ac5, 32'hbeba971b, 32'h3eeb8abf, 32'h3e0a9ada, 32'hbde5e007, 32'hbe1f325e, 32'hbf2ea245, 32'hbed3ae17, 32'hbed6087f, 32'h3ea141fa, 32'hbed0ef58, 32'hbf0f26fa, 32'hbef47265, 32'hbdaf0d62, 32'hbecc5e25, 32'h3daac1ca, 32'h3e53f770, 32'hbecdfb24, 32'hbf158976, 32'hbe7fb1d0, 32'h3e6c2781, 32'hbe026b84, 32'h3e76d330, 32'h3f569124, 32'hbe4b2052, 32'hbf215417, 32'hbeb64fbc, 32'h3ea27ba9, 32'hbd7d8078, 32'h3eaab5df, 32'h3f5c9181, 32'hbec8b20e, 32'hbed528e5, 32'hbed8ce57, 32'hbe83ffc1, 32'hbe12ca22, 32'h3f1a7451, 32'h3f447ab1, 32'hbf09153d, 32'hbf4165ca, 32'hbf207116, 32'hbf059546, 32'h3da9b632, 32'h3ec52774, 32'h3f083d02, 32'hbf9baee6, 32'hbf9fc57d, 32'hbed14d21, 32'hbdd7715a, 32'h3e959824, 32'h3f0748f7, 32'h3f1decea, 32'hbf7839ce, 32'hbf526aae, 32'hbe05fc5f, 32'h3dbf3283, 32'hbdb082bd, 32'hbd2f0a8b, 32'h3ef9a04f, 32'hbf0ce387, 32'hbe6fd3e3, 32'hbe881500, 32'h3d6e035a, 32'h3de8943b, 32'hbcb691ec, 32'h3e4b79c3, 32'h3d89d26e, 32'hbe818460, 32'hbde54390, 32'h3dc15fcc, 32'h3d4828cd, 32'h3caa6298, 32'h3f182573, 32'h3fa91491, 32'h3d2370a0, 32'h3ea9663e, 32'h3f0e3277, 32'hbe011738, 32'hbe9e0be4, 32'hbd93d1a9, 32'hbebfd93b, 32'h3d894c8c, 32'h3e2a34fd, 32'h3e55d095, 32'h3dadb1ab, 32'hbb4c809b, 32'h3f0590dc, 32'h3dbe1c3a, 32'hbe2e064e, 32'hbee37bfd, 32'hbf2d16b7, 32'hbf0a29f7, 32'hbd5da2fe, 32'hbe063250, 32'hbebca124, 32'h3a5b6cd6, 32'hbef87fb3, 32'hbef86f93, 32'hbeed7282, 32'hbe91c4ba, 32'hbe2693f2, 32'h3e2dffa2, 32'hbe5d1090, 32'hbf7054e1, 32'hbefa7869, 32'h3ed45707, 32'hbdd706b4, 32'h3e931e63, 32'h3e06fe8f, 32'h3ee2fd55, 32'hbee54808, 32'hbe9fb639, 32'h3e318b14, 32'h3e447afc, 32'h3d1d5e43, 32'hbbeca9d2, 32'h3f0b50b9, 32'h3d9f97c4, 32'h3f32c86c, 32'h3e506d02, 32'hbd45eb83, 32'hbe49bc24, 32'hbeae2797, 32'hbf089e51, 32'hbead168c, 32'hbe30c061, 32'h3e237d56, 32'h3d668d8b, 32'hbdf22b48, 32'hbe0049ef, 32'hbedf82fc, 32'hbe9c3a94, 32'h3e23db14, 32'h3ed582af, 32'h3ed7c532, 32'h3d41315f, 32'h3eb5d501, 32'hbeb8f0c4, 32'hbeb1072d, 32'hbe452180, 32'h3eaafa59, 32'h3eb210b7, 32'h3e2d3467, 32'hbc3411e0, 32'hbf2851ed, 32'h3e69f9b7, 32'h3e8883cf, 32'h3f0af1a3, 32'h3f512930, 32'h3dc52c39, 32'h3de4b9c3, 32'h3db5f75e, 32'hbe01b675, 32'hbe73b461, 32'h3e9f7bee, 32'h3f114ee3, 32'hbddb3c91, 32'h3cb642f4, 32'hbd8f23f8, 32'h3a807414, 32'h3dac348d, 32'h3eb12c13, 32'h3ebeea7e, 32'hbd817e4c, 32'h3d84c081, 32'hbf270556, 32'h3d5a4fd8, 32'h3e923874, 32'h3f58661c, 32'h3e9f802b, 32'h3ecb2b77, 32'hbd61b59d, 32'hbeaf82a0, 32'hbf673034, 32'hbf19e361, 32'h3d76be78, 32'h3ca759ed, 32'hbe1886ac, 32'hbe6b045f, 32'hbeeafe99, 32'hbf25a2f4, 32'hbe41b8fc, 32'h3c0e8c61, 32'h3eb4c7e2, 32'h3e4ec5de, 32'h3e4e9dc9, 32'h3f0a5ca8, 32'hbeffae7f, 32'hbe457560, 32'hbbdd0b68, 32'h3eace01d, 32'h3ebabeb4, 32'hbdaffd98, 32'hbde53e4f, 32'h3e06a678, 32'hbdd83710, 32'h3e99fb11, 32'h3e1c394e, 32'h3ee64c2a, 32'h3e4da632, 32'h3e939dd4, 32'h3f02353b, 32'hbe18dea5, 32'hbe049697, 32'h3ecc3e53, 32'h3ebc2f92, 32'h3f2841ff, 32'h3f19b192, 32'h3efaf7c4, 32'hbec1fe55, 32'h3e506f43, 32'h3eb4c9b0, 32'h3f241a0f, 32'h3e95e0a2, 32'h3f0ee6b0, 32'h3e360771, 32'hbebdc9c9, 32'hbef802da, 32'h3e731ed0, 32'h3cbb10fb, 32'h3d82e714, 32'hbdb3883a, 32'hbe02c849, 32'hbee3f1a7, 32'hbecd6a9a, 32'h3e18b404, 32'hbe9f9c58, 32'h3c08fd12, 32'h3e0eed68, 32'hbe7821aa, 32'hbd63b2c1, 32'hbf1be7e6, 32'h3ddcd7f8, 32'h3e03c4fd, 32'h3d9dfc5c, 32'h3f410852, 32'h3efe9818, 32'hbd1ec1f6, 32'hbe3c916f, 32'hbe5ff9f0, 32'h3e82eda7, 32'h3e1b5c49, 32'h3d6405fe, 32'h3f0d87d4, 32'h3f412869, 32'hbc9f8d6e, 32'h3f17e4e4, 32'hbf02c509, 32'hbd4e87a8, 32'h3d101660, 32'h3de08274, 32'h3e8e06f0, 32'hbe2f72be, 32'h3df47eb9, 32'h3e0a7fd2, 32'hbe72b77b, 32'h3f130901, 32'h3e977d86, 32'hbe70211a, 32'hbd18dedd, 32'h3e2651c4, 32'h3f3631d4, 32'h3eabfaa6, 32'hbd292843, 32'h3be8f916, 32'hbe284792, 32'hbefcebcd, 32'hbde3490b, 32'hbd391954, 32'hbd0c26fc, 32'h3e78a0db, 32'hbe87de1c, 32'hbe6c8446, 32'hbf3ca3ff, 32'h3e7f772c, 32'h3f2d47f4, 32'h3ed971e2, 32'h3da81e20, 32'h3e147ad7, 32'hbe8b2678, 32'hbf255e76, 32'h3d97492b, 32'h3f5f67c1, 32'h3e73b971, 32'h3ed1a8d6, 32'hbd34c5d1, 32'hbe6422d0, 32'hbec4e713, 32'h3f80651e, 32'h3f755fdd, 32'h3f4c1de2, 32'h3f8aabc2, 32'h3da1cbcf, 32'hbee6c63d, 32'hbf1cc6c0, 32'h3f844b94, 32'h3f7fc20a, 32'h3f9c99bf, 32'h3ed736c2, 32'hbdb154a7, 32'hbe41c039, 32'hbf072581, 32'h3f3d6e59, 32'h3f8b25af, 32'h3f18e496, 32'h3edfea23, 32'h3e08b7c6, 32'hbdab2683, 32'hbefc17eb, 32'h3dc05b39, 32'h3deb4273, 32'h3eb89389, 32'h3ea99ab9, 32'h3d9182f7, 32'hbe7edf2c, 32'hbedc2aa7, 32'h3d32b40b, 32'h3e968049, 32'h3e655965, 32'hbcd08fb9, 32'hbd9f3501, 32'hbdc267d9, 32'hbf33dc0b, 32'h3f61f836, 32'h3f09f405, 32'h3d84ab9a, 32'h3e4ff1c0, 32'h3ef979a5, 32'hbd23c3f3, 32'h3d867a7a, 32'h3eaec8ca, 32'h3f081083, 32'hbd1e74ce, 32'h3e33809b, 32'h3ec3115f, 32'hbf202eca, 32'hbe9280d1, 32'h3e84c5fc, 32'h3e5203da, 32'h3e3b915e, 32'hbbd24204, 32'hbe9ca2ba, 32'h3ea7675e, 32'hbd34494a, 32'hbd33a5cc, 32'h3ee50a6f, 32'hbdca76ee, 32'hbd9c3900, 32'hbec54910, 32'hbe8b3bbe, 32'hbe6bfd56, 32'hbed52ba3, 32'h3f3218ec, 32'h3cb5911d, 32'hbe9467aa, 32'hbe7a2665, 32'hbf46c835, 32'h3d63571d, 32'hbe042aa6, 32'hbdc65c4c, 32'hbf135f44, 32'hbf2a2cdf, 32'hbf10c0d7, 32'hbe95825d, 32'hbe84d91a, 32'h3df38822, 32'hbed322d7, 32'hbf114743, 32'hbf033ad3, 32'h3d5d4b89, 32'h3b543ee5, 32'h3d570a70, 32'h3e766b03, 32'hbe755ba7, 32'hbda7f6d3, 32'hbec9350e, 32'hbd91e85d, 32'h3eb842d0, 32'h3e17dc34, 32'h3d46ed18, 32'h3e16ee16, 32'h3f0e27b0, 32'h3d188dd0, 32'hbde6201c, 32'h3e090d65, 32'hbe4ba0af, 32'hbdec99b8, 32'hbe23b196, 32'h3cc0d397, 32'hbe0a8661, 32'hbf1119cf, 32'h3d760bd6, 32'hbe8b2a0f, 32'hbdbe80bd, 32'hbf04fd89, 32'h3f207f14, 32'hbe9eddb8, 32'h3f328be8, 32'h3ed7a606, 32'h3e886326, 32'h3ebef63c, 32'h3ee957e8, 32'h3e8e1e34, 32'hbebf0ad7, 32'hbed48ab6, 32'h3ebc5d68, 32'hbf0fdfba, 32'hbe4fed43, 32'h3e34acc3, 32'h3e24c3f2, 32'hbebeb9e8, 32'hbf18b8d8, 32'h3e026230, 32'hbe3d6fad, 32'h3e0419f5, 32'hbe2469f8, 32'h3eda4b0f, 32'h3e125a26, 32'h3e253985, 32'h3f04fdbd, 32'h3ebe6083, 32'h3ea5c433, 32'h3e2958ed, 32'hbe880e18, 32'h3e228a56, 32'hbdc4fbfe, 32'hbcd908e2, 32'h3f1064f2, 32'hbe196d68, 32'h3e5c3451, 32'h3f43bf8b, 32'h3e5777b7, 32'hbe8cdf0c, 32'hbe7e76ed, 32'hbda1aa96, 32'hbf38d90f, 32'hbec661c8, 32'h3ebe5c7e, 32'h3e0bd24b, 32'h3da4f7de, 32'h3e071235, 32'hbed64a34, 32'hbebcdfa8, 32'hbdb30bce, 32'h3dc30a1e, 32'h3d602a0d, 32'h3d29e4a7, 32'h3ecf7be9, 32'h3c0bc0bf, 32'hbe96f5f5, 32'h3e87a5c8, 32'h3ed08315, 32'h3e94e976, 32'hbe83813f, 32'h3af06836, 32'hbcf236a3, 32'hbf7710d1, 32'hbeb5b3d4, 32'h3da22636, 32'h3eb89584, 32'hbd9b19f6, 32'hbbe1b377, 32'h3e55a78c, 32'h3db9720e, 32'h3cd45186, 32'h3e788cb3, 32'h3f143c91, 32'h3e652e76, 32'hbd510924, 32'h3f26ba13, 32'hbe235781, 32'hbd9495bf, 32'h3d83ec3c, 32'hbf4827cb, 32'h3f095dbe, 32'h3f21a831, 32'h3e4e1766, 32'h3e4eb873, 32'h3ef64889, 32'h3e93a647, 32'h3df311a3, 32'hbe059155, 32'h3ef9bbcf, 32'h3e9b5472, 32'h3de3fe88, 32'h3f3f44e1, 32'h3eb7ced8, 32'hbdeb21e1, 32'hbeece9ba, 32'h3c4b2bc4, 32'h3f844119, 32'h3fa614dc, 32'h3f003a79, 32'hbd2c1a5d, 32'hbeb0a41c, 32'h3d68aaa5, 32'hbe0959af, 32'h3c9f294a, 32'h3edf9e8a, 32'hbdc82146, 32'hbeb83aa3, 32'h3d2b6050, 32'hbd992bcd, 32'h3e9278c4, 32'hbb4cf218, 32'hbf15aa59, 32'hbc124d73, 32'hbd837256, 32'h3e5917c3, 32'h3dc2b71b, 32'h3f43eb17, 32'hbe5b8338, 32'hbf3ef8e8, 32'hbee8f5b6, 32'h3e8b5533, 32'h3c8a99b2, 32'hbe24f9ee, 32'h3de9470f, 32'hbf342274, 32'hbeda818f, 32'hbf4ed1f5, 32'hbee0c282, 32'hbe1e30d9, 32'hbf33c3ae, 32'hbf0de052, 32'h3e2863cd, 32'h3e6011cc, 32'h3ee1ade2, 32'h3ec70412, 32'hbdc2bfe8, 32'h3e18ee9c, 32'h3e6e5e18, 32'hbd47c910, 32'h3d8bb11a, 32'h3eba5356, 32'hbe9f7935, 32'hbec065f1, 32'hbe7882ec, 32'h3e925d1c, 32'hbe023301, 32'h3eff3119, 32'h3da35a4b, 32'h3eb19b67, 32'hbe713243, 32'h3cfd88f1, 32'hbe7b361f, 32'hbdf3f700, 32'h3d58a0fd, 32'hbec09f87, 32'h3ebaaa32, 32'h3edd7a1d, 32'hbe28a88b, 32'h3ee21ea0, 32'h3e147e1b, 32'hbe1110f0, 32'hbef0fdce, 32'hbf016bfb, 32'h3d5eba6e, 32'h3e2994e4, 32'h3d99e3fd, 32'hbe157648, 32'hbe80cb5f, 32'hbef2f88c, 32'hbd1ac191, 32'h3d79e0e0, 32'h3f0ee882, 32'h3b972fc3, 32'hbe466a18, 32'hbdd2e7fb, 32'h3efd4afd, 32'h3f0a4b9f, 32'h3ef9b02a, 32'h3f031d24, 32'h3f3e8f21, 32'h3efcaecd, 32'h3eab4814, 32'h3d7cb6ac, 32'h3e473fcf, 32'hbdbf5b8d, 32'hbeb8c50d, 32'hbdde6d76, 32'h3f033b77, 32'h3e658b35, 32'h3e6758fc, 32'h3f1ec341, 32'hbf12fb9d, 32'hbf2e1a4a, 32'hbf020cab, 32'h3f0236e3, 32'h3ea6e78c, 32'hbdcda188, 32'hbe79040d, 32'hbd6de126, 32'hbf1f558e, 32'hbf68a820, 32'h3f67ca28, 32'h3e1be6a3, 32'h3ecafbe1, 32'hbe3096f6, 32'hbe39436d, 32'hbef60885, 32'hbea63541, 32'h3f894c43, 32'h3ee80348, 32'hbee5d10d, 32'hbe9ea23b, 32'hbf7ac335, 32'hbe504073, 32'hbed5346e, 32'h3f0a2b8c, 32'hbe20d7f8, 32'hbeb88aa6, 32'hbe60a010, 32'hbea47b4c, 32'hbf006d84, 32'hbda3f67a, 32'h3cc95f6c, 32'hbed1061f, 32'hbcd3d62c, 32'h3f0d0e5e, 32'h3da10c47, 32'hbe32591f, 32'hbede36d4, 32'h3f3aea1f, 32'h3f20d148, 32'h3c00d0a0, 32'hbe73d4a1, 32'hbe015c54, 32'hbd81bbad, 32'h3d2dbd41, 32'h3f1f982a, 32'h3dac6bc7, 32'hbf05947d, 32'hbf487913, 32'hbf1c7746, 32'hbf7e301d, 32'hbf3fcc83, 32'h3cb5be40, 32'h3e920b02, 32'h3e11aa40, 32'hbd4c8f07, 32'hbf2b0c99, 32'hbf1bd341, 32'hbe147484, 32'hbd7c461c, 32'hbeb836b6, 32'hbeb6a9f7, 32'hbeb440b9, 32'hbf3e9108, 32'hbf2056fe, 32'hbe375c13, 32'hbed7bb9d, 32'h3e9f81d3, 32'h3ec7304d, 32'hbdc4c52b, 32'hbf1f0c74, 32'hbebfaaa8, 32'hbee4751b, 32'hbea6b9de, 32'h3f150cb8, 32'h3ef18a02, 32'hbe4f7643, 32'hbeda2152, 32'hb9f39b9b, 32'hbdb338ec, 32'h3e52c7f3, 32'h3f616e30, 32'h3f442268, 32'h3e89d233, 32'h3e8abd67, 32'h3e85b1f0, 32'h3ddc1b32, 32'h3ef3a1d1, 32'h3f16feb2, 32'h3ea2000e, 32'hbd6dbebe, 32'h3e65ed1d, 32'h3f2fb4b5, 32'h3e239311, 32'h3f2b2048, 32'h3dd86b52, 32'hbc7413f3, 32'hbeb6f0f5, 32'h3e7d901e, 32'h3f1cdca1, 32'h3ed275af, 32'hbe71ace9, 32'hbe46715e, 32'h3d913ff6, 32'hbdc3d760, 32'h3d9b5603, 32'hbdd2f271, 32'h3e3c7d67, 32'hbde83e3a, 32'hbeca811b, 32'h3ec12df0, 32'h3d930554, 32'h3f0383ff, 32'hbe8a08df, 32'hbf197962, 32'hbb9dda5b, 32'h3d83aeba, 32'h3f079f99, 32'h3ea03039, 32'hbf23c75c, 32'hbf13820c, 32'hbf868011, 32'hbe1794a5, 32'h3ddee146, 32'h3ed2aa31, 32'hbe54b9f9, 32'hbf412984, 32'hbf1a4f72, 32'hbe7131f3, 32'hbef0f484, 32'hbea70e15, 32'hbe2fca5a, 32'hbf0f2ee1, 32'hbe5fb719, 32'h3b174f11, 32'hbeaf7a2c, 32'hbf1324a2, 32'hbf4bd376, 32'h3f1e9e6a, 32'h3dc012f1, 32'h3ee9e1c5, 32'hbd873522, 32'hbeb4bdd9, 32'h3ee7527e, 32'h3e8330c5, 32'h3e8397d2, 32'hbe0fda06, 32'h3ee50927, 32'hbe06eee2, 32'hbebeb7a5, 32'h3e67f339, 32'h3e78cbcb, 32'h3db3ab25, 32'h3e88111b, 32'h3e482fab, 32'h3e3a72a3, 32'hbe08f620, 32'h3e3d06a6, 32'h3eb9725d, 32'h3f16cf44, 32'hbf009c95, 32'h3e3eda9a, 32'hbf1669ff, 32'hbef27bb7, 32'hbe765f10, 32'h3e675a61, 32'hbedd5a5f, 32'hbe9806df, 32'h3ed5bcb6, 32'hbdfe8c97, 32'hbed7ce8e, 32'h3e6eabfe, 32'h3df80ec2, 32'hbeb40e17, 32'hbe3eb3fd, 32'hbdad59ea, 32'h3e3e8b44, 32'hbeefcc30, 32'hbf0e9f6a, 32'hbeb215e3, 32'hbde293ed, 32'hbeaea9ba, 32'hbe8fd9b7, 32'hbe9a3ad6, 32'hbf1226dc, 32'hbf0ec4ca, 32'h3da858af, 32'h3d5999f4, 32'h3f63acc4, 32'hbe103699, 32'hbd3f2029, 32'hbeb83c95, 32'hbf402156, 32'hbec80513, 32'hbe937289, 32'hbd572790, 32'hbe78d8e5, 32'h3e642146, 32'h3da183c8, 32'hbe848a47, 32'h3e186696, 32'h3f0f4f0b, 32'hbe6879b3, 32'hbed3af8d, 32'h3e119f07, 32'h3ecb9015, 32'h3e64c282, 32'hbef30545, 32'hbebbe098, 32'hbe3dd9bd, 32'hbc73544d, 32'h3f550ff7, 32'h3f0a666a, 32'h3ed58f30, 32'hbf0a2b03, 32'hbecd3caf, 32'h3dc866a4, 32'hbccfe4d5, 32'h3e01f8a6, 32'h3e8c43c7, 32'h3df76ebd, 32'h3d52073c, 32'hbf2b8240, 32'hbd543541, 32'h3e8bf87e, 32'h3d8c82b6, 32'h3edd4b43, 32'h3eb5bf7d, 32'hbf1bb1ff, 32'hbf165bc1, 32'h3d86cfe6, 32'h3e92e04c, 32'hbe4885d6, 32'hbda7baa3, 32'hbf7b7baa, 32'hbf48d829, 32'hbf0649d4, 32'h3d85dd4c, 32'h3ebe3c40, 32'h3c329274, 32'hbead6af5, 32'h3dd557f9, 32'h3ef0f556, 32'hbde2eb83, 32'h3f08a2a7, 32'hbdbc4e21, 32'hbd9d2368, 32'hbea6ede5, 32'h3df0c425, 32'h3df84abb, 32'hbd0c70c8, 32'hbdd216f5, 32'h3cbfb138, 32'hbd1c14ff, 32'hbd8406b9, 32'hbf3401fd, 32'hbf1bbb97, 32'h3e9df599, 32'hbe830251, 32'hbefea280, 32'h3ba8b87f, 32'hbf04c77c, 32'h3f1f3066, 32'h3da7af28, 32'hbe52a117, 32'hbe00fd1e, 32'h3db8ed08, 32'h3d5c8ece, 32'hbe8a3e9e, 32'hbeeba05b, 32'h3eaf81f8, 32'hbf8a9338, 32'h3eb59350, 32'h3f0189b9, 32'h3ef92bb8, 32'hbe37ebd4, 32'hbef66a40, 32'h3e4e4d0c, 32'h3e5546e8, 32'h3c373309, 32'h3d9463d0, 32'h3e0f2d50, 32'hbee876b4, 32'h3eb44024, 32'h3dd47905, 32'h3e720599, 32'hbe193b21, 32'hbcc5e998, 32'h3f8f0c8d, 32'h3edda2c7, 32'h3e6940fc, 32'hbe743a8c, 32'hbf4241f7, 32'hbe9f40f4, 32'hbdbe8e11, 32'h3e3cd70a, 32'hbe8fa19f, 32'h3e5f58ba, 32'hbd0f0073, 32'hbedcb110, 32'h3ee0910f, 32'h3ea5dc21, 32'h3c384a9d, 32'hbdf2a8ee, 32'h3e7edc3d, 32'h3edf3dc3, 32'hbebc68e0, 32'hbf1c0b20, 32'h3ee70a2f, 32'h3ecd2802, 32'hbebea660, 32'h3e918ac1, 32'hbf44d79e, 32'hbf3e18db, 32'hbf66b050, 32'hbd5e5ce1, 32'hbeaf25ac, 32'hbe214756, 32'h3eb2b15e, 32'hbe36be75, 32'hbf288d8b, 32'h3e293107, 32'hbed98927, 32'h3e291b6d, 32'hbc185397, 32'h3ed5813b, 32'h3e20eee8, 32'hbe7fe381, 32'hbe9712b2, 32'hbf0e1a02, 32'h3e46e806, 32'h3e85bf79, 32'h3ece388f, 32'h3e309993, 32'hbd10faa3, 32'hbecd4c43, 32'h3c6aa098, 32'h3ebe19b9, 32'h3f1140cb, 32'hbdf9b716, 32'h3cef97ba, 32'h3e4c6ad0, 32'hbe107a90, 32'h3d656882, 32'hbe47b183, 32'hbf067daa, 32'hbeba94cf, 32'h3e885c56, 32'h3f1921ad, 32'h3f264df4, 32'h3f0fd5bb, 32'h3ea1cc0e, 32'hbf05d88a, 32'hbefff13c, 32'hbe77b537, 32'h3f0a15af, 32'h3f1442fb, 32'hbe1f48c8, 32'hbe68bca5, 32'hbded580a, 32'hbe507ea2, 32'hbe4ed140, 32'hbe79977b, 32'h3cebc2ce, 32'hbf09c112, 32'hbf4ed431, 32'hbf532b0d, 32'hbee78527, 32'hbe9ec31a, 32'h3f0fec3b, 32'h3f2a811f, 32'h3efb8f50, 32'hbe2cd180, 32'hbf5da3a3, 32'hbe6f242c, 32'hbd761f84, 32'h3ec0a233, 32'h3f2671c1, 32'h3eb81ae4, 32'h3bc44330, 32'hbe536d52, 32'hbee1fbc4, 32'hbeb66a9f, 32'hbe1a482d, 32'hbca77c88, 32'hbe868aac, 32'h3dcc1752, 32'hbe68c3ca, 32'h3f821ebd, 32'hbf00da31, 32'hbe46d287, 32'h3e99c53e, 32'hbe87ef49, 32'hbe6b6506, 32'h3edcf9f9, 32'hbd98999a, 32'hbf1199ce, 32'h3e2b4861, 32'h3e43ea8d, 32'h3c2cc3ec, 32'hbd9bc1ae, 32'h3f066f39, 32'hbb5b4205, 32'hbe8cb8e7, 32'hbedaf796, 32'hbf242d23, 32'hbc900836, 32'hbdc10198, 32'hbe095947, 32'hbf09f0a8, 32'h3e9b95f3, 32'hbe02ab28, 32'h3e39d421, 32'h3c63eced, 32'hbebad9cb, 32'hbe55a603, 32'hbe8df75b, 32'h3e9cbae3, 32'hbdba4176, 32'hbe131c01, 32'h3ebba56e, 32'hbf3d6a34, 32'hbebabfd8, 32'h3ed26e67, 32'h3eecd52d, 32'h3e489bca, 32'h3dcf85be, 32'h3d56fd88, 32'hbf0dc2e0, 32'h3e1916e3, 32'h3e88357c, 32'h3e971615, 32'h3e5540fd, 32'hbdb2cfe3, 32'hbee8ef05, 32'hbe4afd10, 32'hbe806e51, 32'h3dd88199, 32'h3f304cc6, 32'h3e845e18, 32'hbd00e79a, 32'h3e9fdbb7, 32'hbeb13332, 32'hbb8196a2, 32'hbeddf83c, 32'hbf10507f, 32'h3d929223, 32'h3e461bf8, 32'h3ec1c72d, 32'hbd6fd48a, 32'h3dd1393b, 32'h3ebaf292, 32'hbe2f456d, 32'hbe100219, 32'h3e292a8e, 32'hbf0451de, 32'hbf4c6b48, 32'hbe967e9a, 32'hbe20e8a6, 32'h3ecb7da6, 32'h3ec20bc3, 32'hbecd5d7b, 32'hbec09627, 32'hbecb98c9, 32'hbe475d28, 32'h3e878f78, 32'h3e9cd138, 32'hbcf57f63, 32'hbf539a4f, 32'hbf24ba80, 32'h3e8ba28f, 32'h3e68f6ed, 32'h3ebd07ba, 32'hbdc766e6, 32'hbe1fba66, 32'hbf0ec117, 32'hbdc5483e, 32'h3ed2454c, 32'h3ed49147, 32'h3e7f03ae, 32'hbd834cc6, 32'hbec1cb98, 32'h3e1cb232, 32'h3f3d3c42, 32'h3d2a8b55, 32'hbe8bfc43, 32'hbe95914a, 32'hbed0cc38, 32'hbed472ee, 32'hbe8139a2, 32'hbf055db8, 32'hbef3b240, 32'h3e4c6431, 32'h3ee471ef, 32'h3f25a664, 32'h3e957c9b, 32'hbeb7be92, 32'hbe93d471, 32'hbebbc231, 32'h3e46df45, 32'hbcddae2f, 32'h3e1f0693, 32'h3e80f289, 32'hbf059b57, 32'hbe96c740, 32'hbf6ff1bb, 32'h3dd50930, 32'h3eca5eaf, 32'h3e0cd587, 32'hbd33eaa7, 32'hbddd79c9, 32'hbedb6d38, 32'hbe078478, 32'h3e9eaa45, 32'h3f417b3c, 32'h3f0b43a3, 32'h3f448cb0, 32'hbd0941ea, 32'h3cecebf2, 32'hbed27188, 32'h3f6e0a3b, 32'h3e0d1958, 32'h3f5ea2bd, 32'h3f3c8dc3, 32'hbdec96ea, 32'hbefe96a6, 32'h3e133a10, 32'h3e4ece07, 32'h3ec77a48, 32'h3f805f77, 32'h3ed1e6d0, 32'hbeb33bda, 32'hbeb5ba95, 32'hbdb52389, 32'h3cbd82b2, 32'h3eb49b90, 32'h3f140ee7, 32'hbe3d5d8a};

    localparam integer positions[0:49][1:2] = '{
        '{0,1850},
        '{50,1888},
        '{100,1926},
        '{150,1964},
        '{200,2002},
        '{250,0},
        '{300,0},
        '{350,0},
        '{400,0},
        '{450,0},
        '{500,0},
        '{550,0},
        '{600,0},
        '{650,0},
        '{700,0},
        '{750,0},
        '{800,0},
        '{850,0},
        '{900,0},
        '{950,0},
        '{1000,0},
        '{1050,0},
        '{1100,0},
        '{1150,0},
        '{1200,0},
        '{1250,0},
        '{1300,0},
        '{1350,0},
        '{1400,0},
        '{1450,0},
        '{1500,0},
        '{1550,0},
        '{1600,0},
        '{1650,0},
        '{1700,0},
        '{1750,0},
        '{1800,0},
        '{1850,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0},
        '{0,0}
    };

endpackage