--
--##################################
--#extended for different bit width# -> choose bit width for sigmoid 
--##################################
--
-- megafunction wizard: %ROM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: sigmoid_IP.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2020  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and any partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details, at
--https://fpgasoftware.intel.com/eula.
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
--
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;
--
ENTITY sigmoid_IP IS
	PORT
	(
--		
--choose bit width for sigmoid 
		--address : IN STD_LOGIC_VECTOR ( 2 DOWNTO 0); -- 3 Bit
		--address : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0); -- 4 Bit		
		--address : IN STD_LOGIC_VECTOR ( 4 DOWNTO 0); -- 5 Bit
		--address : IN STD_LOGIC_VECTOR ( 5 DOWNTO 0); -- 6 Bit
		--address : IN STD_LOGIC_VECTOR ( 6 DOWNTO 0); -- 7 Bit
		--address : IN STD_LOGIC_VECTOR ( 7 DOWNTO 0); -- 8 Bit
		--address : IN STD_LOGIC_VECTOR ( 8 DOWNTO 0); -- 9 Bit
		--address : IN STD_LOGIC_VECTOR ( 9 DOWNTO 0); --10 Bit		
		--address : IN STD_LOGIC_VECTOR (10 DOWNTO 0); --11 Bit
		address : IN STD_LOGIC_VECTOR (11 DOWNTO 0); --12 Bit	
--
		clock		: IN STD_LOGIC  := '1';
		q		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END sigmoid_IP;
--
ARCHITECTURE SYN OF sigmoid_ip IS
--
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (7 DOWNTO 0);
--
BEGIN
	q    <= sub_wire0(7 DOWNTO 0);
--
	altsyncram_component : altsyncram
	GENERIC MAP (
		address_aclr_a => "NONE",
		clock_enable_input_a => "BYPASS",
		clock_enable_output_a => "BYPASS",
--		
--choose bit width for sigmoid
		--init_file => "sigmoid_3_bit.mif",  -- 3 Bit
		--init_file => "sigmoid_4_bit.mif",  -- 4 Bit
		--init_file => "sigmoid_5_bit.mif",  -- 5 Bit
		--init_file => "sigmoid_6_bit.mif",  -- 6 Bit
		--init_file => "sigmoid_7_bit.mif",  -- 7 Bit
		--init_file => "sigmoid_8_bit.mif",  -- 8 Bit
		--init_file => "sigmoid_9_bit.mif",  -- 9 Bit
		--init_file => "sigmoid_10_bit.mif", --10 Bit
		--init_file => "sigmoid_11_bit.mif", --11 Bit
		init_file => "sigmoid_values.mif", --12 Bit
--
		intended_device_family => "Cyclone IV E",
		lpm_hint => "ENABLE_RUNTIME_MOD=NO",
		lpm_type => "altsyncram",
--
--choose bit width for sigmoid
		--numwords_a =>    8, -- 3 Bit
		--numwords_a =>   16, -- 4 Bit
		--numwords_a =>   32, -- 5 Bit
		--numwords_a =>   64, -- 6 Bit
		--numwords_a =>  128, -- 7 Bit
		--numwords_a =>  256, -- 8 Bit
		--numwords_a =>  512, -- 9 Bit		
		--numwords_a => 1024, --10 Bit
		--numwords_a => 2048, --11 Bit
		numwords_a => 4096, --12 Bit 
--		
		operation_mode => "ROM",
		outdata_aclr_a => "NONE",
		outdata_reg_a => "CLOCK0",
--		
--choose bit width for sigmoid		
		--widthad_a =>  3, -- 3 Bit		
		--widthad_a =>  4, -- 4 Bit
		--widthad_a =>  5, -- 5 Bit
		--widthad_a =>  6, -- 6 Bit
		--widthad_a =>  7, -- 7 Bit
		--widthad_a =>  8, -- 8 Bit
		--widthad_a =>  9, -- 9 Bit
		--widthad_a => 10, --10 Bit
		--widthad_a => 11, --11 Bit
		widthad_a => 12, --12 Bit
--
		width_a => 8,
		width_byteena_a => 1
	)
	PORT MAP (
		address_a => address,
		clock0 => clock,
		q_a => sub_wire0
	);
--
END SYN;
--
-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
-- Retrieval info: PRIVATE: AclrAddr NUMERIC "0"
-- Retrieval info: PRIVATE: AclrByte NUMERIC "0"
-- Retrieval info: PRIVATE: AclrOutput NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
-- Retrieval info: PRIVATE: BlankMemory NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "0"
-- Retrieval info: PRIVATE: Clken NUMERIC "0"
-- Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
-- Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
-- Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
-- Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
-- Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
-- Retrieval info: PRIVATE: MIFfilename STRING "sigmoid_12_bit.mif"
-- Retrieval info: PRIVATE: NUMWORDS_A NUMERIC "4096"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: RegAddr NUMERIC "1"
-- Retrieval info: PRIVATE: RegOutput NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: SingleClock NUMERIC "1"
-- Retrieval info: PRIVATE: UseDQRAM NUMERIC "0"
-- Retrieval info: PRIVATE: WidthAddr NUMERIC "12"
-- Retrieval info: PRIVATE: WidthData NUMERIC "8"
-- Retrieval info: PRIVATE: rden NUMERIC "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: ADDRESS_ACLR_A STRING "NONE"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "BYPASS"
-- Retrieval info: CONSTANT: INIT_FILE STRING "sigmoid_12_bit.mif"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: LPM_HINT STRING "ENABLE_RUNTIME_MOD=NO"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
-- Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "4096"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "ROM"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
-- Retrieval info: CONSTANT: OUTDATA_REG_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "12"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
-- Retrieval info: USED_PORT: address 0 0 12 0 INPUT NODEFVAL "address[11..0]"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT VCC "clock"
-- Retrieval info: USED_PORT: q 0 0 8 0 OUTPUT NODEFVAL "q[7..0]"
-- Retrieval info: CONNECT: @address_a 0 0 12 0 address 0 0 12 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: q 0 0 8 0 @q_a 0 0 8 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL sigmoid_IP.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sigmoid_IP.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sigmoid_IP.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sigmoid_IP.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sigmoid_IP_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
